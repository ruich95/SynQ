module rv32i (
    input wire clk,
    input wire [0:0] w_0,
    input wire [31:0] w_1,
    input wire [31:0] w_2,
    output wire [0:0] w_1616,
    output wire [31:0] w_1617,
    output wire [31:0] w_1618,
    output wire [31:0] w_1619);

  wire [31:0] w_3;
  wire [31:0] w_4;
  wire [31:0] w_5;
  wire [31:0] w_6;
  wire [31:0] w_7;
  wire [31:0] w_8;
  wire [31:0] w_9;
  wire [31:0] w_10;
  wire [31:0] w_11;
  wire [31:0] w_12;
  wire [31:0] w_13;
  wire [31:0] w_14;
  wire [31:0] w_15;
  wire [31:0] w_16;
  wire [31:0] w_17;
  wire [31:0] w_18;
  wire [31:0] w_19;
  wire [31:0] w_20;
  wire [31:0] w_21;
  wire [31:0] w_22;
  wire [31:0] w_23;
  wire [31:0] w_24;
  wire [31:0] w_25;
  wire [31:0] w_26;
  wire [31:0] w_27;
  wire [31:0] w_28;
  wire [31:0] w_29;
  wire [31:0] w_30;
  wire [31:0] w_31;
  wire [31:0] w_32;
  wire [31:0] w_33;
  wire [31:0] w_34;
  wire [31:0] w_264;
  wire [31:0] w_265;
  wire [31:0] w_266;
  wire [31:0] w_267;
  wire [31:0] w_268;
  wire [31:0] w_269;
  wire [31:0] w_270;
  wire [31:0] w_271;
  wire [31:0] w_272;
  wire [31:0] w_273;
  wire [31:0] w_274;
  wire [31:0] w_275;
  wire [31:0] w_276;
  wire [31:0] w_277;
  wire [31:0] w_278;
  wire [31:0] w_279;
  wire [31:0] w_280;
  wire [31:0] w_281;
  wire [31:0] w_282;
  wire [31:0] w_283;
  wire [31:0] w_284;
  wire [31:0] w_285;
  wire [31:0] w_286;
  wire [31:0] w_287;
  wire [31:0] w_288;
  wire [31:0] w_289;
  wire [31:0] w_290;
  wire [31:0] w_291;
  wire [31:0] w_292;
  wire [31:0] w_293;
  wire [31:0] w_294;
  wire [31:0] w_295;
  wire [31:0] w_389;
  wire [31:0] w_390;
  wire [31:0] w_391;
  wire [31:0] w_392;
  wire [31:0] w_393;
  wire [31:0] w_394;
  wire [31:0] w_395;
  wire [31:0] w_396;
  wire [31:0] w_397;
  wire [31:0] w_398;
  wire [31:0] w_399;
  wire [31:0] w_400;
  wire [31:0] w_401;
  wire [31:0] w_402;
  wire [31:0] w_403;
  wire [31:0] w_404;
  wire [31:0] w_405;
  wire [31:0] w_406;
  wire [31:0] w_407;
  wire [31:0] w_408;
  wire [31:0] w_409;
  wire [31:0] w_410;
  wire [31:0] w_411;
  wire [31:0] w_412;
  wire [31:0] w_413;
  wire [31:0] w_414;
  wire [31:0] w_415;
  wire [31:0] w_416;
  wire [31:0] w_417;
  wire [31:0] w_418;
  wire [31:0] w_419;
  wire [31:0] w_420;
  wire [31:0] w_421;
  wire [4:0] w_229;
  wire [31:0] w_230;
  wire [31:0] w_231;
  wire [31:0] w_232;
  wire [31:0] w_233;
  wire [31:0] w_234;
  wire [31:0] w_235;
  wire [31:0] w_236;
  wire [31:0] w_237;
  wire [31:0] w_238;
  wire [31:0] w_239;
  wire [31:0] w_240;
  wire [31:0] w_241;
  wire [31:0] w_242;
  wire [31:0] w_243;
  wire [31:0] w_244;
  wire [31:0] w_245;
  wire [31:0] w_246;
  wire [31:0] w_247;
  wire [31:0] w_248;
  wire [31:0] w_249;
  wire [31:0] w_250;
  wire [31:0] w_251;
  wire [31:0] w_252;
  wire [31:0] w_253;
  wire [31:0] w_254;
  wire [31:0] w_255;
  wire [31:0] w_256;
  wire [31:0] w_257;
  wire [31:0] w_258;
  wire [31:0] w_259;
  wire [31:0] w_260;
  wire [31:0] w_261;
  wire [31:0] w_193;
  wire [4:0] w_194;
  wire [31:0] w_195;
  wire [31:0] w_196;
  wire [31:0] w_197;
  wire [31:0] w_198;
  wire [31:0] w_199;
  wire [31:0] w_200;
  wire [31:0] w_201;
  wire [31:0] w_202;
  wire [31:0] w_203;
  wire [31:0] w_204;
  wire [31:0] w_205;
  wire [31:0] w_206;
  wire [31:0] w_207;
  wire [31:0] w_208;
  wire [31:0] w_209;
  wire [31:0] w_210;
  wire [31:0] w_211;
  wire [31:0] w_212;
  wire [31:0] w_213;
  wire [31:0] w_214;
  wire [31:0] w_215;
  wire [31:0] w_216;
  wire [31:0] w_217;
  wire [31:0] w_218;
  wire [31:0] w_219;
  wire [31:0] w_220;
  wire [31:0] w_221;
  wire [31:0] w_222;
  wire [31:0] w_223;
  wire [31:0] w_224;
  wire [31:0] w_225;
  wire [31:0] w_226;
  wire [31:0] w_159;
  wire [31:0] w_160;
  wire [31:0] w_161;
  wire [31:0] w_162;
  wire [31:0] w_163;
  wire [31:0] w_164;
  wire [31:0] w_165;
  wire [31:0] w_166;
  wire [31:0] w_167;
  wire [31:0] w_168;
  wire [31:0] w_169;
  wire [31:0] w_170;
  wire [31:0] w_171;
  wire [31:0] w_172;
  wire [31:0] w_173;
  wire [31:0] w_174;
  wire [31:0] w_175;
  wire [31:0] w_176;
  wire [31:0] w_177;
  wire [31:0] w_178;
  wire [31:0] w_179;
  wire [31:0] w_180;
  wire [31:0] w_181;
  wire [31:0] w_182;
  wire [31:0] w_183;
  wire [31:0] w_184;
  wire [31:0] w_185;
  wire [31:0] w_186;
  wire [31:0] w_187;
  wire [31:0] w_188;
  wire [31:0] w_189;
  wire [31:0] w_190;
  wire [31:0] w_191;
  wire [32:0] w_640;
  wire [32:0] w_645;
  wire [32:0] w_650;
  wire [32:0] w_689;
  wire [32:0] w_692;
  wire [0:0] w_657;
  wire [0:0] w_658;
  wire [0:0] w_659;
  wire [32:0] w_696;
  wire [32:0] w_834;
  wire [32:0] w_842;
  wire [32:0] w_887;
  wire [32:0] w_892;
  wire [32:0] w_895;
  wire [9:0] w_879;
  wire [31:0] w_471;
  wire [31:0] w_882;
  wire [32:0] w_1323;
  wire [31:0] w_594;
  wire [31:0] w_457;
  wire [31:0] w_458;
  wire [0:0] w_465;
  wire [0:0] w_466;
  wire [4:0] w_467;
  wire [31:0] w_468;
  wire [31:0] w_469;
  wire [2:0] w_470;
  wire [0:0] w_1356;
  wire [0:0] w_1357;
  wire [4:0] w_1358;
  wire [31:0] w_1359;
  wire [31:0] w_1360;
  wire [2:0] w_1361;
  wire [0:0] w_1343;
  wire [0:0] w_1344;
  wire [4:0] w_1345;
  wire [31:0] w_1346;
  wire [31:0] w_1347;
  wire [2:0] w_1348;
  wire [0:0] w_1337;
  wire [31:0] w_1338;
  wire [31:0] w_1339;
  wire [31:0] w_1340;
  wire [4:0] w_1341;
  wire [31:0] w_1342;
  wire [0:0] w_1362;
  wire [0:0] w_1363;
  wire [4:0] w_1364;
  wire [31:0] w_1365;
  wire [31:0] w_1366;
  wire [2:0] w_1367;
  wire [0:0] w_599;
  wire [31:0] w_633;
  wire [31:0] w_704;
  wire [4:0] w_727;
  wire [31:0] w_1297;
  wire [0:0] w_1306;
  wire [0:0] w_1312;
  wire [4:0] w_1319;
  wire [31:0] w_1321;
  wire [31:0] w_1326;
  wire [2:0] w_1329;
  wire [0:0] w_1330;
  wire [0:0] w_1331;
  wire [4:0] w_1332;
  wire [31:0] w_1333;
  wire [31:0] w_1334;
  wire [2:0] w_1335;
  wire [0:0] w_459;
  wire [0:0] w_460;
  wire [4:0] w_461;
  wire [31:0] w_462;
  wire [31:0] w_463;
  wire [2:0] w_464;
  wire [31:0] w_228;
  wire [31:0] w_423;
  wire [31:0] w_1453;
  wire [31:0] w_1455;
  wire [31:0] w_1457;
  wire [31:0] w_1459;
  wire [31:0] w_1461;
  wire [31:0] w_1463;
  wire [31:0] w_1465;
  wire [31:0] w_1467;
  wire [31:0] w_1469;
  wire [31:0] w_1471;
  wire [31:0] w_1473;
  wire [31:0] w_1475;
  wire [31:0] w_1477;
  wire [31:0] w_1479;
  wire [31:0] w_1481;
  wire [31:0] w_1483;
  wire [31:0] w_1485;
  wire [31:0] w_1487;
  wire [31:0] w_1489;
  wire [31:0] w_1491;
  wire [31:0] w_1493;
  wire [31:0] w_1495;
  wire [31:0] w_1497;
  wire [31:0] w_1499;
  wire [31:0] w_1501;
  wire [31:0] w_1503;
  wire [31:0] w_1505;
  wire [31:0] w_1507;
  wire [31:0] w_1509;
  wire [31:0] w_1511;
  wire [31:0] w_1513;
  wire [31:0] w_1451;
  wire [31:0] w_1388;
  wire [31:0] w_1389;
  wire [31:0] w_1390;
  wire [31:0] w_1391;
  wire [31:0] w_1392;
  wire [31:0] w_1393;
  wire [31:0] w_1394;
  wire [31:0] w_1395;
  wire [31:0] w_1396;
  wire [31:0] w_1397;
  wire [31:0] w_1398;
  wire [31:0] w_1399;
  wire [31:0] w_1400;
  wire [31:0] w_1401;
  wire [31:0] w_1402;
  wire [31:0] w_1403;
  wire [31:0] w_1404;
  wire [31:0] w_1405;
  wire [31:0] w_1406;
  wire [31:0] w_1407;
  wire [31:0] w_1408;
  wire [31:0] w_1409;
  wire [31:0] w_1410;
  wire [31:0] w_1411;
  wire [31:0] w_1412;
  wire [31:0] w_1413;
  wire [31:0] w_1414;
  wire [31:0] w_1415;
  wire [31:0] w_1416;
  wire [31:0] w_1417;
  wire [31:0] w_1418;
  wire [31:0] w_1419;
  wire [31:0] w_1547;
  wire [31:0] w_1548;
  wire [31:0] w_1549;
  wire [31:0] w_1550;
  wire [31:0] w_1551;
  wire [31:0] w_1552;
  wire [31:0] w_1553;
  wire [31:0] w_1554;
  wire [31:0] w_1555;
  wire [31:0] w_1556;
  wire [31:0] w_1557;
  wire [31:0] w_1558;
  wire [31:0] w_1559;
  wire [31:0] w_1560;
  wire [31:0] w_1561;
  wire [31:0] w_1562;
  wire [31:0] w_1563;
  wire [31:0] w_1564;
  wire [31:0] w_1565;
  wire [31:0] w_1566;
  wire [31:0] w_1567;
  wire [31:0] w_1568;
  wire [31:0] w_1569;
  wire [31:0] w_1570;
  wire [31:0] w_1571;
  wire [31:0] w_1572;
  wire [31:0] w_1573;
  wire [31:0] w_1574;
  wire [31:0] w_1575;
  wire [31:0] w_1576;
  wire [31:0] w_1577;
  wire [31:0] w_1578;
  wire [0:0] w_1612;
  wire [31:0] w_1613;
  wire [31:0] w_1614;
  wire [31:0] w_1615;
  wire [0:0] w_1382;
  wire [31:0] w_1383;
  wire [31:0] w_1384;
  wire [31:0] w_1385;
  wire [0:0] w_1369;
  wire [31:0] w_1370;
  wire [31:0] w_1371;
  wire [31:0] w_1372;
  wire [4:0] w_1373;
  wire [31:0] w_1374;
  wire [31:0] w_424;
  wire [31:0] w_425;
  wire [31:0] w_426;
  wire [31:0] w_427;
  wire [31:0] w_428;
  wire [31:0] w_429;
  wire [31:0] w_430;
  wire [31:0] w_431;
  wire [31:0] w_432;
  wire [31:0] w_433;
  wire [31:0] w_434;
  wire [31:0] w_435;
  wire [31:0] w_436;
  wire [31:0] w_437;
  wire [31:0] w_438;
  wire [31:0] w_439;
  wire [31:0] w_440;
  wire [31:0] w_441;
  wire [31:0] w_442;
  wire [31:0] w_443;
  wire [31:0] w_444;
  wire [31:0] w_445;
  wire [31:0] w_446;
  wire [31:0] w_447;
  wire [31:0] w_448;
  wire [31:0] w_449;
  wire [31:0] w_450;
  wire [31:0] w_451;
  wire [31:0] w_452;
  wire [31:0] w_453;
  wire [31:0] w_454;
  wire [31:0] w_455;
  wire [0:0] w_1375;
  wire [0:0] w_1376;
  wire [4:0] w_1377;
  wire [31:0] w_1378;
  wire [31:0] w_1379;
  wire [2:0] w_1380;
  wire [31:0] w_35;
  wire [31:0] w_36;
  wire [31:0] w_37;
  wire [31:0] w_38;
  wire [31:0] w_39;
  wire [31:0] w_40;
  wire [31:0] w_41;
  wire [31:0] w_42;
  wire [31:0] w_43;
  wire [31:0] w_44;
  wire [31:0] w_45;
  wire [31:0] w_46;
  wire [31:0] w_47;
  wire [31:0] w_48;
  wire [31:0] w_49;
  wire [31:0] w_50;
  wire [31:0] w_51;
  wire [31:0] w_52;
  wire [31:0] w_53;
  wire [31:0] w_54;
  wire [31:0] w_55;
  wire [31:0] w_56;
  wire [31:0] w_57;
  wire [31:0] w_58;
  wire [31:0] w_59;
  wire [31:0] w_60;
  wire [31:0] w_61;
  wire [31:0] w_62;
  wire [31:0] w_63;
  wire [31:0] w_64;
  wire [31:0] w_65;
  wire [31:0] w_66;
  wire [31:0] w_296;
  wire [31:0] w_297;
  wire [31:0] w_298;
  wire [31:0] w_299;
  wire [31:0] w_300;
  wire [31:0] w_301;
  wire [31:0] w_302;
  wire [31:0] w_303;
  wire [31:0] w_304;
  wire [31:0] w_305;
  wire [31:0] w_306;
  wire [31:0] w_307;
  wire [31:0] w_308;
  wire [31:0] w_309;
  wire [31:0] w_310;
  wire [31:0] w_311;
  wire [31:0] w_312;
  wire [31:0] w_313;
  wire [31:0] w_314;
  wire [31:0] w_315;
  wire [31:0] w_316;
  wire [31:0] w_317;
  wire [31:0] w_318;
  wire [31:0] w_319;
  wire [31:0] w_320;
  wire [31:0] w_321;
  wire [31:0] w_322;
  wire [31:0] w_323;
  wire [31:0] w_324;
  wire [31:0] w_325;
  wire [31:0] w_326;
  wire [31:0] w_327;
  wire [4:0] w_263;
  wire [32:0] w_641;
  wire [32:0] w_646;
  wire [32:0] w_651;
  wire [32:0] w_690;
  wire [32:0] w_693;
  wire [0:0] w_660;
  wire [0:0] w_661;
  wire [0:0] w_662;
  wire [32:0] w_697;
  wire [32:0] w_835;
  wire [32:0] w_843;
  wire [32:0] w_888;
  wire [32:0] w_893;
  wire [32:0] w_896;
  wire [9:0] w_883;
  wire [31:0] w_884;
  wire [31:0] w_885;
  wire [32:0] w_1324;
  wire [31:0] w_595;
  wire [31:0] w_472;
  wire [0:0] w_473;
  wire [0:0] w_474;
  wire [4:0] w_475;
  wire [31:0] w_476;
  wire [31:0] w_477;
  wire [2:0] w_478;
  wire [0:0] w_1349;
  wire [0:0] w_1350;
  wire [4:0] w_1351;
  wire [31:0] w_1352;
  wire [31:0] w_1353;
  wire [2:0] w_1354;
  wire [31:0] w_1420;
  wire [31:0] w_1421;
  wire [31:0] w_1422;
  wire [31:0] w_1423;
  wire [31:0] w_1424;
  wire [31:0] w_1425;
  wire [31:0] w_1426;
  wire [31:0] w_1427;
  wire [31:0] w_1428;
  wire [31:0] w_1429;
  wire [31:0] w_1430;
  wire [31:0] w_1431;
  wire [31:0] w_1432;
  wire [31:0] w_1433;
  wire [31:0] w_1434;
  wire [31:0] w_1435;
  wire [31:0] w_1436;
  wire [31:0] w_1437;
  wire [31:0] w_1438;
  wire [31:0] w_1439;
  wire [31:0] w_1440;
  wire [31:0] w_1441;
  wire [31:0] w_1442;
  wire [31:0] w_1443;
  wire [31:0] w_1444;
  wire [31:0] w_1445;
  wire [31:0] w_1446;
  wire [31:0] w_1447;
  wire [31:0] w_1448;
  wire [31:0] w_1449;
  wire [31:0] w_1450;
  wire [31:0] w_1514;
  wire [31:0] w_1515;
  wire [31:0] w_1516;
  wire [31:0] w_1517;
  wire [31:0] w_1518;
  wire [31:0] w_1519;
  wire [31:0] w_1520;
  wire [31:0] w_1521;
  wire [31:0] w_1522;
  wire [31:0] w_1523;
  wire [31:0] w_1524;
  wire [31:0] w_1525;
  wire [31:0] w_1526;
  wire [31:0] w_1527;
  wire [31:0] w_1528;
  wire [31:0] w_1529;
  wire [31:0] w_1530;
  wire [31:0] w_1531;
  wire [31:0] w_1532;
  wire [31:0] w_1533;
  wire [31:0] w_1534;
  wire [31:0] w_1535;
  wire [31:0] w_1536;
  wire [31:0] w_1537;
  wire [31:0] w_1538;
  wire [31:0] w_1539;
  wire [31:0] w_1540;
  wire [31:0] w_1541;
  wire [31:0] w_1542;
  wire [31:0] w_1543;
  wire [31:0] w_1544;
  wire [31:0] w_1545;
  wire [31:0] w_1579;
  wire [31:0] w_1580;
  wire [31:0] w_1581;
  wire [31:0] w_1582;
  wire [31:0] w_1583;
  wire [31:0] w_1584;
  wire [31:0] w_1585;
  wire [31:0] w_1586;
  wire [31:0] w_1587;
  wire [31:0] w_1588;
  wire [31:0] w_1589;
  wire [31:0] w_1590;
  wire [31:0] w_1591;
  wire [31:0] w_1592;
  wire [31:0] w_1593;
  wire [31:0] w_1594;
  wire [31:0] w_1595;
  wire [31:0] w_1596;
  wire [31:0] w_1597;
  wire [31:0] w_1598;
  wire [31:0] w_1599;
  wire [31:0] w_1600;
  wire [31:0] w_1601;
  wire [31:0] w_1602;
  wire [31:0] w_1603;
  wire [31:0] w_1604;
  wire [31:0] w_1605;
  wire [31:0] w_1606;
  wire [31:0] w_1607;
  wire [31:0] w_1608;
  wire [31:0] w_1609;
  wire [31:0] w_1610;
  wire [4:0] w_1386;
  wire [31:0] w_1387;
  wire [0:0] w_1620;
  wire [0:0] w_1621;
  wire [4:0] w_1622;
  wire [31:0] w_1623;
  wire [31:0] w_1624;
  wire [2:0] w_1625;
  wire [4:0] w_67;
  wire [0:0] w_68;
  wire [4:0] w_69;
  wire [0:0] w_70;
  wire [4:0] w_71;
  wire [0:0] w_72;
  wire [4:0] w_73;
  wire [0:0] w_74;
  wire [4:0] w_75;
  wire [0:0] w_76;
  wire [4:0] w_77;
  wire [0:0] w_78;
  wire [4:0] w_79;
  wire [0:0] w_80;
  wire [4:0] w_81;
  wire [0:0] w_82;
  wire [4:0] w_83;
  wire [0:0] w_84;
  wire [4:0] w_85;
  wire [0:0] w_86;
  wire [4:0] w_87;
  wire [0:0] w_88;
  wire [4:0] w_89;
  wire [0:0] w_90;
  wire [4:0] w_91;
  wire [0:0] w_92;
  wire [4:0] w_93;
  wire [0:0] w_94;
  wire [4:0] w_95;
  wire [0:0] w_96;
  wire [4:0] w_97;
  wire [0:0] w_98;
  wire [4:0] w_99;
  wire [0:0] w_100;
  wire [4:0] w_101;
  wire [0:0] w_102;
  wire [4:0] w_103;
  wire [0:0] w_104;
  wire [4:0] w_105;
  wire [0:0] w_106;
  wire [4:0] w_107;
  wire [0:0] w_108;
  wire [4:0] w_109;
  wire [0:0] w_110;
  wire [4:0] w_111;
  wire [0:0] w_112;
  wire [4:0] w_113;
  wire [0:0] w_114;
  wire [4:0] w_115;
  wire [0:0] w_116;
  wire [4:0] w_117;
  wire [0:0] w_118;
  wire [4:0] w_119;
  wire [0:0] w_120;
  wire [4:0] w_121;
  wire [0:0] w_122;
  wire [4:0] w_123;
  wire [0:0] w_124;
  wire [4:0] w_125;
  wire [0:0] w_126;
  wire [4:0] w_127;
  wire [0:0] w_128;
  wire [31:0] w_129;
  wire [31:0] w_130;
  wire [31:0] w_131;
  wire [31:0] w_132;
  wire [31:0] w_133;
  wire [31:0] w_134;
  wire [31:0] w_135;
  wire [31:0] w_136;
  wire [31:0] w_137;
  wire [31:0] w_138;
  wire [31:0] w_139;
  wire [31:0] w_140;
  wire [31:0] w_141;
  wire [31:0] w_142;
  wire [31:0] w_143;
  wire [31:0] w_144;
  wire [31:0] w_145;
  wire [31:0] w_146;
  wire [31:0] w_147;
  wire [31:0] w_148;
  wire [31:0] w_149;
  wire [31:0] w_150;
  wire [31:0] w_151;
  wire [31:0] w_152;
  wire [31:0] w_153;
  wire [31:0] w_154;
  wire [31:0] w_155;
  wire [31:0] w_156;
  wire [31:0] w_157;
  wire [31:0] w_158;
  wire [0:0] w_328;
  wire [0:0] w_329;
  wire [0:0] w_330;
  wire [0:0] w_331;
  wire [0:0] w_332;
  wire [0:0] w_333;
  wire [0:0] w_334;
  wire [0:0] w_335;
  wire [0:0] w_336;
  wire [0:0] w_337;
  wire [0:0] w_338;
  wire [0:0] w_339;
  wire [0:0] w_340;
  wire [0:0] w_341;
  wire [0:0] w_342;
  wire [0:0] w_343;
  wire [0:0] w_344;
  wire [0:0] w_345;
  wire [0:0] w_346;
  wire [0:0] w_347;
  wire [0:0] w_348;
  wire [0:0] w_349;
  wire [0:0] w_350;
  wire [0:0] w_351;
  wire [0:0] w_352;
  wire [0:0] w_353;
  wire [0:0] w_354;
  wire [0:0] w_355;
  wire [0:0] w_356;
  wire [0:0] w_357;
  wire [0:0] w_358;
  wire [31:0] w_359;
  wire [31:0] w_360;
  wire [31:0] w_361;
  wire [31:0] w_362;
  wire [31:0] w_363;
  wire [31:0] w_364;
  wire [31:0] w_365;
  wire [31:0] w_366;
  wire [31:0] w_367;
  wire [31:0] w_368;
  wire [31:0] w_369;
  wire [31:0] w_370;
  wire [31:0] w_371;
  wire [31:0] w_372;
  wire [31:0] w_373;
  wire [31:0] w_374;
  wire [31:0] w_375;
  wire [31:0] w_376;
  wire [31:0] w_377;
  wire [31:0] w_378;
  wire [31:0] w_379;
  wire [31:0] w_380;
  wire [31:0] w_381;
  wire [31:0] w_382;
  wire [31:0] w_383;
  wire [31:0] w_384;
  wire [31:0] w_385;
  wire [31:0] w_386;
  wire [31:0] w_387;
  wire [31:0] w_388;
  wire [6:0] w_479;
  wire [0:0] w_480;
  wire [6:0] w_481;
  wire [0:0] w_482;
  wire [6:0] w_483;
  wire [0:0] w_484;
  wire [0:0] w_485;
  wire [0:0] w_486;
  wire [6:0] w_487;
  wire [4:0] w_488;
  wire [11:0] w_489;
  wire [0:0] w_490;
  wire [19:0] w_491;
  wire [19:0] w_492;
  wire [6:0] w_493;
  wire [4:0] w_494;
  wire [11:0] w_495;
  wire [31:0] w_496;
  wire [6:0] w_497;
  wire [0:0] w_498;
  wire [6:0] w_499;
  wire [4:0] w_500;
  wire [11:0] w_501;
  wire [0:0] w_502;
  wire [19:0] w_503;
  wire [19:0] w_504;
  wire [6:0] w_505;
  wire [4:0] w_506;
  wire [11:0] w_507;
  wire [31:0] w_508;
  wire [6:0] w_509;
  wire [0:0] w_510;
  wire [6:0] w_511;
  wire [0:0] w_512;
  wire [4:0] w_513;
  wire [0:0] w_514;
  wire [1:0] w_515;
  wire [6:0] w_516;
  wire [5:0] w_517;
  wire [4:0] w_518;
  wire [4:0] w_519;
  wire [4:0] w_520;
  wire [10:0] w_521;
  wire [12:0] w_522;
  wire [0:0] w_523;
  wire [18:0] w_524;
  wire [18:0] w_525;
  wire [6:0] w_526;
  wire [0:0] w_527;
  wire [4:0] w_528;
  wire [0:0] w_529;
  wire [1:0] w_530;
  wire [6:0] w_531;
  wire [5:0] w_532;
  wire [4:0] w_533;
  wire [4:0] w_534;
  wire [4:0] w_535;
  wire [10:0] w_536;
  wire [12:0] w_537;
  wire [31:0] w_538;
  wire [6:0] w_539;
  wire [0:0] w_540;
  wire [6:0] w_541;
  wire [0:0] w_542;
  wire [0:0] w_543;
  wire [6:0] w_544;
  wire [4:0] w_545;
  wire [11:0] w_546;
  wire [4:0] w_547;
  wire [2:0] w_548;
  wire [7:0] w_549;
  wire [19:0] w_550;
  wire [31:0] w_551;
  wire [6:0] w_552;
  wire [0:0] w_553;
  wire [6:0] w_554;
  wire [0:0] w_555;
  wire [4:0] w_556;
  wire [2:0] w_557;
  wire [7:0] w_558;
  wire [8:0] w_559;
  wire [4:0] w_560;
  wire [0:0] w_561;
  wire [6:0] w_562;
  wire [5:0] w_563;
  wire [4:0] w_564;
  wire [4:0] w_565;
  wire [4:0] w_566;
  wire [10:0] w_567;
  wire [11:0] w_568;
  wire [20:0] w_569;
  wire [0:0] w_570;
  wire [10:0] w_571;
  wire [10:0] w_572;
  wire [6:0] w_573;
  wire [0:0] w_574;
  wire [4:0] w_575;
  wire [2:0] w_576;
  wire [7:0] w_577;
  wire [8:0] w_578;
  wire [4:0] w_579;
  wire [0:0] w_580;
  wire [6:0] w_581;
  wire [5:0] w_582;
  wire [4:0] w_583;
  wire [4:0] w_584;
  wire [4:0] w_585;
  wire [10:0] w_586;
  wire [11:0] w_587;
  wire [20:0] w_588;
  wire [31:0] w_589;
  wire [31:0] w_590;
  wire [31:0] w_591;
  wire [31:0] w_592;
  wire [31:0] w_593;
  wire [0:0] w_596;
  wire [0:0] w_597;
  wire [0:0] w_598;
  wire [0:0] w_600;
  wire [6:0] w_601;
  wire [4:0] w_602;
  wire [11:0] w_603;
  wire [4:0] w_604;
  wire [2:0] w_605;
  wire [7:0] w_606;
  wire [19:0] w_607;
  wire [4:0] w_608;
  wire [6:0] w_609;
  wire [11:0] w_610;
  wire [31:0] w_611;
  wire [15:0] w_612;
  wire [15:0] w_613;
  wire [31:0] w_614;
  wire [0:0] w_615;
  wire [6:0] w_616;
  wire [4:0] w_617;
  wire [11:0] w_618;
  wire [4:0] w_619;
  wire [2:0] w_620;
  wire [7:0] w_621;
  wire [19:0] w_622;
  wire [4:0] w_623;
  wire [6:0] w_624;
  wire [11:0] w_625;
  wire [31:0] w_626;
  wire [23:0] w_627;
  wire [7:0] w_628;
  wire [31:0] w_629;
  wire [31:0] w_630;
  wire [31:0] w_631;
  wire [31:0] w_632;
  wire [0:0] w_634;
  wire [6:0] w_635;
  wire [0:0] w_636;
  wire [6:0] w_637;
  wire [0:0] w_638;
  wire [0:0] w_639;
  wire [31:0] w_642;
  wire [6:0] w_643;
  wire [0:0] w_644;
  wire [31:0] w_647;
  wire [6:0] w_648;
  wire [0:0] w_649;
  wire [31:0] w_652;
  wire [31:0] w_653;
  wire [31:0] w_654;
  wire [6:0] w_655;
  wire [0:0] w_656;
  wire [2:0] w_663;
  wire [0:0] w_664;
  wire [0:0] w_665;
  wire [2:0] w_666;
  wire [0:0] w_667;
  wire [0:0] w_668;
  wire [0:0] w_669;
  wire [0:0] w_670;
  wire [2:0] w_671;
  wire [0:0] w_672;
  wire [0:0] w_673;
  wire [2:0] w_674;
  wire [0:0] w_675;
  wire [0:0] w_676;
  wire [0:0] w_677;
  wire [0:0] w_678;
  wire [2:0] w_679;
  wire [0:0] w_680;
  wire [0:0] w_681;
  wire [2:0] w_682;
  wire [0:0] w_683;
  wire [0:0] w_684;
  wire [0:0] w_685;
  wire [0:0] w_686;
  wire [0:0] w_687;
  wire [0:0] w_688;
  wire [31:0] w_691;
  wire [31:0] w_694;
  wire [31:0] w_695;
  wire [31:0] w_698;
  wire [31:0] w_699;
  wire [31:0] w_700;
  wire [31:0] w_701;
  wire [31:0] w_702;
  wire [31:0] w_703;
  wire [0:0] w_705;
  wire [4:0] w_706;
  wire [6:0] w_707;
  wire [0:0] w_708;
  wire [6:0] w_709;
  wire [0:0] w_710;
  wire [0:0] w_711;
  wire [6:0] w_712;
  wire [0:0] w_713;
  wire [6:0] w_714;
  wire [0:0] w_715;
  wire [0:0] w_716;
  wire [0:0] w_717;
  wire [6:0] w_718;
  wire [0:0] w_719;
  wire [6:0] w_720;
  wire [0:0] w_721;
  wire [0:0] w_722;
  wire [0:0] w_723;
  wire [4:0] w_724;
  wire [4:0] w_725;
  wire [4:0] w_726;
  wire [0:0] w_728;
  wire [6:0] w_729;
  wire [4:0] w_730;
  wire [11:0] w_731;
  wire [4:0] w_732;
  wire [2:0] w_733;
  wire [7:0] w_734;
  wire [19:0] w_735;
  wire [4:0] w_736;
  wire [6:0] w_737;
  wire [11:0] w_738;
  wire [31:0] w_739;
  wire [15:0] w_740;
  wire [0:0] w_741;
  wire [15:0] w_742;
  wire [15:0] w_743;
  wire [6:0] w_744;
  wire [4:0] w_745;
  wire [11:0] w_746;
  wire [4:0] w_747;
  wire [2:0] w_748;
  wire [7:0] w_749;
  wire [19:0] w_750;
  wire [4:0] w_751;
  wire [6:0] w_752;
  wire [11:0] w_753;
  wire [31:0] w_754;
  wire [15:0] w_755;
  wire [31:0] w_756;
  wire [0:0] w_757;
  wire [6:0] w_758;
  wire [4:0] w_759;
  wire [11:0] w_760;
  wire [4:0] w_761;
  wire [2:0] w_762;
  wire [7:0] w_763;
  wire [19:0] w_764;
  wire [4:0] w_765;
  wire [6:0] w_766;
  wire [11:0] w_767;
  wire [31:0] w_768;
  wire [7:0] w_769;
  wire [0:0] w_770;
  wire [23:0] w_771;
  wire [23:0] w_772;
  wire [6:0] w_773;
  wire [4:0] w_774;
  wire [11:0] w_775;
  wire [4:0] w_776;
  wire [2:0] w_777;
  wire [7:0] w_778;
  wire [19:0] w_779;
  wire [4:0] w_780;
  wire [6:0] w_781;
  wire [11:0] w_782;
  wire [31:0] w_783;
  wire [7:0] w_784;
  wire [31:0] w_785;
  wire [0:0] w_786;
  wire [6:0] w_787;
  wire [4:0] w_788;
  wire [11:0] w_789;
  wire [4:0] w_790;
  wire [2:0] w_791;
  wire [7:0] w_792;
  wire [19:0] w_793;
  wire [4:0] w_794;
  wire [6:0] w_795;
  wire [11:0] w_796;
  wire [31:0] w_797;
  wire [15:0] w_798;
  wire [31:0] w_799;
  wire [0:0] w_800;
  wire [6:0] w_801;
  wire [4:0] w_802;
  wire [11:0] w_803;
  wire [4:0] w_804;
  wire [2:0] w_805;
  wire [7:0] w_806;
  wire [19:0] w_807;
  wire [4:0] w_808;
  wire [6:0] w_809;
  wire [11:0] w_810;
  wire [31:0] w_811;
  wire [7:0] w_812;
  wire [31:0] w_813;
  wire [6:0] w_814;
  wire [4:0] w_815;
  wire [11:0] w_816;
  wire [4:0] w_817;
  wire [2:0] w_818;
  wire [7:0] w_819;
  wire [19:0] w_820;
  wire [4:0] w_821;
  wire [6:0] w_822;
  wire [11:0] w_823;
  wire [31:0] w_824;
  wire [31:0] w_825;
  wire [31:0] w_826;
  wire [31:0] w_827;
  wire [31:0] w_828;
  wire [31:0] w_829;
  wire [6:0] w_830;
  wire [0:0] w_831;
  wire [6:0] w_832;
  wire [0:0] w_833;
  wire [31:0] w_836;
  wire [6:0] w_837;
  wire [0:0] w_838;
  wire [6:0] w_839;
  wire [0:0] w_840;
  wire [0:0] w_841;
  wire [31:0] w_844;
  wire [6:0] w_845;
  wire [0:0] w_846;
  wire [6:0] w_847;
  wire [0:0] w_848;
  wire [0:0] w_849;
  wire [2:0] w_850;
  wire [0:0] w_851;
  wire [6:0] w_852;
  wire [0:0] w_853;
  wire [6:0] w_854;
  wire [0:0] w_855;
  wire [9:0] w_856;
  wire [9:0] w_857;
  wire [2:0] w_858;
  wire [0:0] w_859;
  wire [2:0] w_860;
  wire [0:0] w_861;
  wire [2:0] w_862;
  wire [0:0] w_863;
  wire [2:0] w_864;
  wire [0:0] w_865;
  wire [2:0] w_866;
  wire [0:0] w_867;
  wire [6:0] w_868;
  wire [0:0] w_869;
  wire [9:0] w_870;
  wire [2:0] w_871;
  wire [0:0] w_872;
  wire [9:0] w_873;
  wire [9:0] w_874;
  wire [9:0] w_875;
  wire [9:0] w_876;
  wire [9:0] w_877;
  wire [9:0] w_878;
  wire [6:0] w_880;
  wire [0:0] w_881;
  wire [0:0] w_886;
  wire [31:0] w_889;
  wire [0:0] w_890;
  wire [31:0] w_891;
  wire [31:0] w_894;
  wire [31:0] w_897;
  wire [0:0] w_898;
  wire [0:0] w_899;
  wire [31:0] w_900;
  wire [0:0] w_901;
  wire [0:0] w_902;
  wire [31:0] w_903;
  wire [0:0] w_904;
  wire [31:0] w_905;
  wire [0:0] w_906;
  wire [4:0] w_907;
  wire [0:0] w_908;
  wire [31:0] w_909;
  wire [4:0] w_910;
  wire [0:0] w_911;
  wire [31:0] w_912;
  wire [4:0] w_913;
  wire [0:0] w_914;
  wire [31:0] w_915;
  wire [4:0] w_916;
  wire [0:0] w_917;
  wire [31:0] w_918;
  wire [4:0] w_919;
  wire [0:0] w_920;
  wire [31:0] w_921;
  wire [4:0] w_922;
  wire [0:0] w_923;
  wire [31:0] w_924;
  wire [4:0] w_925;
  wire [0:0] w_926;
  wire [31:0] w_927;
  wire [4:0] w_928;
  wire [0:0] w_929;
  wire [31:0] w_930;
  wire [4:0] w_931;
  wire [0:0] w_932;
  wire [31:0] w_933;
  wire [4:0] w_934;
  wire [0:0] w_935;
  wire [31:0] w_936;
  wire [4:0] w_937;
  wire [0:0] w_938;
  wire [31:0] w_939;
  wire [4:0] w_940;
  wire [0:0] w_941;
  wire [31:0] w_942;
  wire [4:0] w_943;
  wire [0:0] w_944;
  wire [31:0] w_945;
  wire [4:0] w_946;
  wire [0:0] w_947;
  wire [31:0] w_948;
  wire [4:0] w_949;
  wire [0:0] w_950;
  wire [31:0] w_951;
  wire [4:0] w_952;
  wire [0:0] w_953;
  wire [31:0] w_954;
  wire [4:0] w_955;
  wire [0:0] w_956;
  wire [31:0] w_957;
  wire [4:0] w_958;
  wire [0:0] w_959;
  wire [31:0] w_960;
  wire [4:0] w_961;
  wire [0:0] w_962;
  wire [31:0] w_963;
  wire [4:0] w_964;
  wire [0:0] w_965;
  wire [31:0] w_966;
  wire [4:0] w_967;
  wire [0:0] w_968;
  wire [31:0] w_969;
  wire [4:0] w_970;
  wire [0:0] w_971;
  wire [31:0] w_972;
  wire [4:0] w_973;
  wire [0:0] w_974;
  wire [31:0] w_975;
  wire [4:0] w_976;
  wire [0:0] w_977;
  wire [31:0] w_978;
  wire [4:0] w_979;
  wire [0:0] w_980;
  wire [31:0] w_981;
  wire [4:0] w_982;
  wire [0:0] w_983;
  wire [31:0] w_984;
  wire [4:0] w_985;
  wire [0:0] w_986;
  wire [31:0] w_987;
  wire [4:0] w_988;
  wire [0:0] w_989;
  wire [31:0] w_990;
  wire [4:0] w_991;
  wire [0:0] w_992;
  wire [31:0] w_993;
  wire [4:0] w_994;
  wire [0:0] w_995;
  wire [31:0] w_996;
  wire [4:0] w_997;
  wire [0:0] w_998;
  wire [31:0] w_999;
  wire [31:0] w_1000;
  wire [31:0] w_1001;
  wire [31:0] w_1002;
  wire [31:0] w_1003;
  wire [31:0] w_1004;
  wire [31:0] w_1005;
  wire [31:0] w_1006;
  wire [31:0] w_1007;
  wire [31:0] w_1008;
  wire [31:0] w_1009;
  wire [31:0] w_1010;
  wire [31:0] w_1011;
  wire [31:0] w_1012;
  wire [31:0] w_1013;
  wire [31:0] w_1014;
  wire [31:0] w_1015;
  wire [31:0] w_1016;
  wire [31:0] w_1017;
  wire [31:0] w_1018;
  wire [31:0] w_1019;
  wire [31:0] w_1020;
  wire [31:0] w_1021;
  wire [31:0] w_1022;
  wire [31:0] w_1023;
  wire [31:0] w_1024;
  wire [31:0] w_1025;
  wire [31:0] w_1026;
  wire [31:0] w_1027;
  wire [31:0] w_1028;
  wire [31:0] w_1029;
  wire [31:0] w_1030;
  wire [0:0] w_1031;
  wire [4:0] w_1032;
  wire [0:0] w_1033;
  wire [31:0] w_1034;
  wire [4:0] w_1035;
  wire [0:0] w_1036;
  wire [31:0] w_1037;
  wire [4:0] w_1038;
  wire [0:0] w_1039;
  wire [31:0] w_1040;
  wire [4:0] w_1041;
  wire [0:0] w_1042;
  wire [31:0] w_1043;
  wire [4:0] w_1044;
  wire [0:0] w_1045;
  wire [31:0] w_1046;
  wire [4:0] w_1047;
  wire [0:0] w_1048;
  wire [31:0] w_1049;
  wire [4:0] w_1050;
  wire [0:0] w_1051;
  wire [31:0] w_1052;
  wire [4:0] w_1053;
  wire [0:0] w_1054;
  wire [31:0] w_1055;
  wire [4:0] w_1056;
  wire [0:0] w_1057;
  wire [31:0] w_1058;
  wire [4:0] w_1059;
  wire [0:0] w_1060;
  wire [31:0] w_1061;
  wire [4:0] w_1062;
  wire [0:0] w_1063;
  wire [31:0] w_1064;
  wire [4:0] w_1065;
  wire [0:0] w_1066;
  wire [31:0] w_1067;
  wire [4:0] w_1068;
  wire [0:0] w_1069;
  wire [31:0] w_1070;
  wire [4:0] w_1071;
  wire [0:0] w_1072;
  wire [31:0] w_1073;
  wire [4:0] w_1074;
  wire [0:0] w_1075;
  wire [31:0] w_1076;
  wire [4:0] w_1077;
  wire [0:0] w_1078;
  wire [31:0] w_1079;
  wire [4:0] w_1080;
  wire [0:0] w_1081;
  wire [31:0] w_1082;
  wire [4:0] w_1083;
  wire [0:0] w_1084;
  wire [31:0] w_1085;
  wire [4:0] w_1086;
  wire [0:0] w_1087;
  wire [31:0] w_1088;
  wire [4:0] w_1089;
  wire [0:0] w_1090;
  wire [31:0] w_1091;
  wire [4:0] w_1092;
  wire [0:0] w_1093;
  wire [31:0] w_1094;
  wire [4:0] w_1095;
  wire [0:0] w_1096;
  wire [31:0] w_1097;
  wire [4:0] w_1098;
  wire [0:0] w_1099;
  wire [31:0] w_1100;
  wire [4:0] w_1101;
  wire [0:0] w_1102;
  wire [31:0] w_1103;
  wire [4:0] w_1104;
  wire [0:0] w_1105;
  wire [31:0] w_1106;
  wire [4:0] w_1107;
  wire [0:0] w_1108;
  wire [31:0] w_1109;
  wire [4:0] w_1110;
  wire [0:0] w_1111;
  wire [31:0] w_1112;
  wire [4:0] w_1113;
  wire [0:0] w_1114;
  wire [31:0] w_1115;
  wire [4:0] w_1116;
  wire [0:0] w_1117;
  wire [31:0] w_1118;
  wire [4:0] w_1119;
  wire [0:0] w_1120;
  wire [31:0] w_1121;
  wire [4:0] w_1122;
  wire [0:0] w_1123;
  wire [31:0] w_1124;
  wire [31:0] w_1125;
  wire [31:0] w_1126;
  wire [31:0] w_1127;
  wire [31:0] w_1128;
  wire [31:0] w_1129;
  wire [31:0] w_1130;
  wire [31:0] w_1131;
  wire [31:0] w_1132;
  wire [31:0] w_1133;
  wire [31:0] w_1134;
  wire [31:0] w_1135;
  wire [31:0] w_1136;
  wire [31:0] w_1137;
  wire [31:0] w_1138;
  wire [31:0] w_1139;
  wire [31:0] w_1140;
  wire [31:0] w_1141;
  wire [31:0] w_1142;
  wire [31:0] w_1143;
  wire [31:0] w_1144;
  wire [31:0] w_1145;
  wire [31:0] w_1146;
  wire [31:0] w_1147;
  wire [31:0] w_1148;
  wire [31:0] w_1149;
  wire [31:0] w_1150;
  wire [31:0] w_1151;
  wire [31:0] w_1152;
  wire [31:0] w_1153;
  wire [31:0] w_1154;
  wire [31:0] w_1155;
  wire [0:0] w_1156;
  wire [4:0] w_1157;
  wire [0:0] w_1158;
  wire [31:0] w_1159;
  wire [4:0] w_1160;
  wire [0:0] w_1161;
  wire [31:0] w_1162;
  wire [4:0] w_1163;
  wire [0:0] w_1164;
  wire [31:0] w_1165;
  wire [4:0] w_1166;
  wire [0:0] w_1167;
  wire [31:0] w_1168;
  wire [4:0] w_1169;
  wire [0:0] w_1170;
  wire [31:0] w_1171;
  wire [4:0] w_1172;
  wire [0:0] w_1173;
  wire [31:0] w_1174;
  wire [4:0] w_1175;
  wire [0:0] w_1176;
  wire [31:0] w_1177;
  wire [4:0] w_1178;
  wire [0:0] w_1179;
  wire [31:0] w_1180;
  wire [4:0] w_1181;
  wire [0:0] w_1182;
  wire [31:0] w_1183;
  wire [4:0] w_1184;
  wire [0:0] w_1185;
  wire [31:0] w_1186;
  wire [4:0] w_1187;
  wire [0:0] w_1188;
  wire [31:0] w_1189;
  wire [4:0] w_1190;
  wire [0:0] w_1191;
  wire [31:0] w_1192;
  wire [4:0] w_1193;
  wire [0:0] w_1194;
  wire [31:0] w_1195;
  wire [4:0] w_1196;
  wire [0:0] w_1197;
  wire [31:0] w_1198;
  wire [4:0] w_1199;
  wire [0:0] w_1200;
  wire [31:0] w_1201;
  wire [4:0] w_1202;
  wire [0:0] w_1203;
  wire [31:0] w_1204;
  wire [4:0] w_1205;
  wire [0:0] w_1206;
  wire [31:0] w_1207;
  wire [4:0] w_1208;
  wire [0:0] w_1209;
  wire [31:0] w_1210;
  wire [4:0] w_1211;
  wire [0:0] w_1212;
  wire [31:0] w_1213;
  wire [4:0] w_1214;
  wire [0:0] w_1215;
  wire [31:0] w_1216;
  wire [4:0] w_1217;
  wire [0:0] w_1218;
  wire [31:0] w_1219;
  wire [4:0] w_1220;
  wire [0:0] w_1221;
  wire [31:0] w_1222;
  wire [4:0] w_1223;
  wire [0:0] w_1224;
  wire [31:0] w_1225;
  wire [4:0] w_1226;
  wire [0:0] w_1227;
  wire [31:0] w_1228;
  wire [4:0] w_1229;
  wire [0:0] w_1230;
  wire [31:0] w_1231;
  wire [4:0] w_1232;
  wire [0:0] w_1233;
  wire [31:0] w_1234;
  wire [4:0] w_1235;
  wire [0:0] w_1236;
  wire [31:0] w_1237;
  wire [4:0] w_1238;
  wire [0:0] w_1239;
  wire [31:0] w_1240;
  wire [4:0] w_1241;
  wire [0:0] w_1242;
  wire [31:0] w_1243;
  wire [4:0] w_1244;
  wire [0:0] w_1245;
  wire [31:0] w_1246;
  wire [4:0] w_1247;
  wire [0:0] w_1248;
  wire [31:0] w_1249;
  wire [31:0] w_1250;
  wire [31:0] w_1251;
  wire [31:0] w_1252;
  wire [31:0] w_1253;
  wire [31:0] w_1254;
  wire [31:0] w_1255;
  wire [31:0] w_1256;
  wire [31:0] w_1257;
  wire [31:0] w_1258;
  wire [31:0] w_1259;
  wire [31:0] w_1260;
  wire [31:0] w_1261;
  wire [31:0] w_1262;
  wire [31:0] w_1263;
  wire [31:0] w_1264;
  wire [31:0] w_1265;
  wire [31:0] w_1266;
  wire [31:0] w_1267;
  wire [31:0] w_1268;
  wire [31:0] w_1269;
  wire [31:0] w_1270;
  wire [31:0] w_1271;
  wire [31:0] w_1272;
  wire [31:0] w_1273;
  wire [31:0] w_1274;
  wire [31:0] w_1275;
  wire [31:0] w_1276;
  wire [31:0] w_1277;
  wire [31:0] w_1278;
  wire [31:0] w_1279;
  wire [31:0] w_1280;
  wire [0:0] w_1281;
  wire [31:0] w_1282;
  wire [31:0] w_1283;
  wire [31:0] w_1284;
  wire [31:0] w_1285;
  wire [31:0] w_1286;
  wire [31:0] w_1287;
  wire [31:0] w_1288;
  wire [31:0] w_1289;
  wire [31:0] w_1290;
  wire [31:0] w_1291;
  wire [31:0] w_1292;
  wire [31:0] w_1293;
  wire [31:0] w_1294;
  wire [31:0] w_1295;
  wire [31:0] w_1296;
  wire [0:0] w_1298;
  wire [6:0] w_1299;
  wire [0:0] w_1300;
  wire [6:0] w_1301;
  wire [0:0] w_1302;
  wire [0:0] w_1303;
  wire [0:0] w_1304;
  wire [0:0] w_1305;
  wire [0:0] w_1307;
  wire [6:0] w_1308;
  wire [0:0] w_1309;
  wire [0:0] w_1310;
  wire [0:0] w_1311;
  wire [0:0] w_1313;
  wire [6:0] w_1314;
  wire [0:0] w_1315;
  wire [4:0] w_1316;
  wire [4:0] w_1317;
  wire [4:0] w_1318;
  wire [0:0] w_1320;
  wire [0:0] w_1322;
  wire [31:0] w_1325;
  wire [0:0] w_1327;
  wire [2:0] w_1328;
  wire [0:0] w_1452;
  wire [0:0] w_1454;
  wire [0:0] w_1456;
  wire [0:0] w_1458;
  wire [0:0] w_1460;
  wire [0:0] w_1462;
  wire [0:0] w_1464;
  wire [0:0] w_1466;
  wire [0:0] w_1468;
  wire [0:0] w_1470;
  wire [0:0] w_1472;
  wire [0:0] w_1474;
  wire [0:0] w_1476;
  wire [0:0] w_1478;
  wire [0:0] w_1480;
  wire [0:0] w_1482;
  wire [0:0] w_1484;
  wire [0:0] w_1486;
  wire [0:0] w_1488;
  wire [0:0] w_1490;
  wire [0:0] w_1492;
  wire [0:0] w_1494;
  wire [0:0] w_1496;
  wire [0:0] w_1498;
  wire [0:0] w_1500;
  wire [0:0] w_1502;
  wire [0:0] w_1504;
  wire [0:0] w_1506;
  wire [0:0] w_1508;
  wire [0:0] w_1510;
  wire [0:0] w_1512;

  reg [31:0] r_3;
  reg [31:0] r_4;
  reg [31:0] r_5;
  reg [31:0] r_6;
  reg [31:0] r_7;
  reg [31:0] r_8;
  reg [31:0] r_9;
  reg [31:0] r_10;
  reg [31:0] r_11;
  reg [31:0] r_12;
  reg [31:0] r_13;
  reg [31:0] r_14;
  reg [31:0] r_15;
  reg [31:0] r_16;
  reg [31:0] r_17;
  reg [31:0] r_18;
  reg [31:0] r_19;
  reg [31:0] r_20;
  reg [31:0] r_21;
  reg [31:0] r_22;
  reg [31:0] r_23;
  reg [31:0] r_24;
  reg [31:0] r_25;
  reg [31:0] r_26;
  reg [31:0] r_27;
  reg [31:0] r_28;
  reg [31:0] r_29;
  reg [31:0] r_30;
  reg [31:0] r_31;
  reg [31:0] r_32;
  reg [31:0] r_33;
  reg [31:0] r_34;
  reg [0:0] r_459;
  reg [0:0] r_460;
  reg [4:0] r_461;
  reg [31:0] r_462;
  reg [31:0] r_463;
  reg [2:0] r_464;

  assign w_3 = r_3;
  assign w_4 = r_4;
  assign w_5 = r_5;
  assign w_6 = r_6;
  assign w_7 = r_7;
  assign w_8 = r_8;
  assign w_9 = r_9;
  assign w_10 = r_10;
  assign w_11 = r_11;
  assign w_12 = r_12;
  assign w_13 = r_13;
  assign w_14 = r_14;
  assign w_15 = r_15;
  assign w_16 = r_16;
  assign w_17 = r_17;
  assign w_18 = r_18;
  assign w_19 = r_19;
  assign w_20 = r_20;
  assign w_21 = r_21;
  assign w_22 = r_22;
  assign w_23 = r_23;
  assign w_24 = r_24;
  assign w_25 = r_25;
  assign w_26 = r_26;
  assign w_27 = r_27;
  assign w_28 = r_28;
  assign w_29 = r_29;
  assign w_30 = r_30;
  assign w_31 = r_31;
  assign w_32 = r_32;
  assign w_33 = r_33;
  assign w_34 = r_34;
  assign w_459 = r_459;
  assign w_460 = r_460;
  assign w_461 = r_461;
  assign w_462 = r_462;
  assign w_463 = r_463;
  assign w_464 = r_464;

  assign w_35 = w_3;
  assign w_36 = w_4;
  assign w_37 = w_5;
  assign w_38 = w_6;
  assign w_39 = w_7;
  assign w_40 = w_8;
  assign w_41 = w_9;
  assign w_42 = w_10;
  assign w_43 = w_11;
  assign w_44 = w_12;
  assign w_45 = w_13;
  assign w_46 = w_14;
  assign w_47 = w_15;
  assign w_48 = w_16;
  assign w_49 = w_17;
  assign w_50 = w_18;
  assign w_51 = w_19;
  assign w_52 = w_20;
  assign w_53 = w_21;
  assign w_54 = w_22;
  assign w_55 = w_23;
  assign w_56 = w_24;
  assign w_57 = w_25;
  assign w_58 = w_26;
  assign w_59 = w_27;
  assign w_60 = w_28;
  assign w_61 = w_29;
  assign w_62 = w_30;
  assign w_63 = w_31;
  assign w_64 = w_32;
  assign w_65 = w_33;
  assign w_66 = w_34;
  assign w_160 = w_3;
  assign w_161 = w_4;
  assign w_162 = w_5;
  assign w_163 = w_6;
  assign w_164 = w_7;
  assign w_165 = w_8;
  assign w_166 = w_9;
  assign w_167 = w_10;
  assign w_168 = w_11;
  assign w_169 = w_12;
  assign w_170 = w_13;
  assign w_171 = w_14;
  assign w_172 = w_15;
  assign w_173 = w_16;
  assign w_174 = w_17;
  assign w_175 = w_18;
  assign w_176 = w_19;
  assign w_177 = w_20;
  assign w_178 = w_21;
  assign w_179 = w_22;
  assign w_180 = w_23;
  assign w_181 = w_24;
  assign w_182 = w_25;
  assign w_183 = w_26;
  assign w_184 = w_27;
  assign w_185 = w_28;
  assign w_186 = w_29;
  assign w_187 = w_30;
  assign w_188 = w_31;
  assign w_189 = w_32;
  assign w_190 = w_33;
  assign w_191 = w_34;
  assign w_296 = w_264;
  assign w_297 = w_265;
  assign w_298 = w_266;
  assign w_299 = w_267;
  assign w_300 = w_268;
  assign w_301 = w_269;
  assign w_302 = w_270;
  assign w_303 = w_271;
  assign w_304 = w_272;
  assign w_305 = w_273;
  assign w_306 = w_274;
  assign w_307 = w_275;
  assign w_308 = w_276;
  assign w_309 = w_277;
  assign w_310 = w_278;
  assign w_311 = w_279;
  assign w_312 = w_280;
  assign w_313 = w_281;
  assign w_314 = w_282;
  assign w_315 = w_283;
  assign w_316 = w_284;
  assign w_317 = w_285;
  assign w_318 = w_286;
  assign w_319 = w_287;
  assign w_320 = w_288;
  assign w_321 = w_289;
  assign w_322 = w_290;
  assign w_323 = w_291;
  assign w_324 = w_292;
  assign w_325 = w_293;
  assign w_326 = w_294;
  assign w_327 = w_295;
  assign w_390 = w_264;
  assign w_391 = w_265;
  assign w_392 = w_266;
  assign w_393 = w_267;
  assign w_394 = w_268;
  assign w_395 = w_269;
  assign w_396 = w_270;
  assign w_397 = w_271;
  assign w_398 = w_272;
  assign w_399 = w_273;
  assign w_400 = w_274;
  assign w_401 = w_275;
  assign w_402 = w_276;
  assign w_403 = w_277;
  assign w_404 = w_278;
  assign w_405 = w_279;
  assign w_406 = w_280;
  assign w_407 = w_281;
  assign w_408 = w_282;
  assign w_409 = w_283;
  assign w_410 = w_284;
  assign w_411 = w_285;
  assign w_412 = w_286;
  assign w_413 = w_287;
  assign w_414 = w_288;
  assign w_415 = w_289;
  assign w_416 = w_290;
  assign w_417 = w_291;
  assign w_418 = w_292;
  assign w_419 = w_293;
  assign w_420 = w_294;
  assign w_421 = w_295;
  assign w_423 = w_389;
  assign w_424 = w_390;
  assign w_425 = w_391;
  assign w_426 = w_392;
  assign w_427 = w_393;
  assign w_428 = w_394;
  assign w_429 = w_395;
  assign w_430 = w_396;
  assign w_431 = w_397;
  assign w_432 = w_398;
  assign w_433 = w_399;
  assign w_434 = w_400;
  assign w_435 = w_401;
  assign w_436 = w_402;
  assign w_437 = w_403;
  assign w_438 = w_404;
  assign w_439 = w_405;
  assign w_440 = w_406;
  assign w_441 = w_407;
  assign w_442 = w_408;
  assign w_443 = w_409;
  assign w_444 = w_410;
  assign w_445 = w_411;
  assign w_446 = w_412;
  assign w_447 = w_413;
  assign w_448 = w_414;
  assign w_449 = w_415;
  assign w_450 = w_416;
  assign w_451 = w_417;
  assign w_452 = w_418;
  assign w_453 = w_419;
  assign w_454 = w_420;
  assign w_455 = w_421;
  assign w_263 = w_229;
  assign w_264 = w_230;
  assign w_265 = w_231;
  assign w_266 = w_232;
  assign w_267 = w_233;
  assign w_268 = w_234;
  assign w_269 = w_235;
  assign w_270 = w_236;
  assign w_271 = w_237;
  assign w_272 = w_238;
  assign w_273 = w_239;
  assign w_274 = w_240;
  assign w_275 = w_241;
  assign w_276 = w_242;
  assign w_277 = w_243;
  assign w_278 = w_244;
  assign w_279 = w_245;
  assign w_280 = w_246;
  assign w_281 = w_247;
  assign w_282 = w_248;
  assign w_283 = w_249;
  assign w_284 = w_250;
  assign w_285 = w_251;
  assign w_286 = w_252;
  assign w_287 = w_253;
  assign w_288 = w_254;
  assign w_289 = w_255;
  assign w_290 = w_256;
  assign w_291 = w_257;
  assign w_292 = w_258;
  assign w_293 = w_259;
  assign w_294 = w_260;
  assign w_295 = w_261;
  assign w_228 = w_193;
  assign w_229 = w_194;
  assign w_230 = w_195;
  assign w_231 = w_196;
  assign w_232 = w_197;
  assign w_233 = w_198;
  assign w_234 = w_199;
  assign w_235 = w_200;
  assign w_236 = w_201;
  assign w_237 = w_202;
  assign w_238 = w_203;
  assign w_239 = w_204;
  assign w_240 = w_205;
  assign w_241 = w_206;
  assign w_242 = w_207;
  assign w_243 = w_208;
  assign w_244 = w_209;
  assign w_245 = w_210;
  assign w_246 = w_211;
  assign w_247 = w_212;
  assign w_248 = w_213;
  assign w_249 = w_214;
  assign w_250 = w_215;
  assign w_251 = w_216;
  assign w_252 = w_217;
  assign w_253 = w_218;
  assign w_254 = w_219;
  assign w_255 = w_220;
  assign w_256 = w_221;
  assign w_257 = w_222;
  assign w_258 = w_223;
  assign w_259 = w_224;
  assign w_260 = w_225;
  assign w_261 = w_226;
  assign w_193 = w_159;
  assign w_195 = w_160;
  assign w_196 = w_161;
  assign w_197 = w_162;
  assign w_198 = w_163;
  assign w_199 = w_164;
  assign w_200 = w_165;
  assign w_201 = w_166;
  assign w_202 = w_167;
  assign w_203 = w_168;
  assign w_204 = w_169;
  assign w_205 = w_170;
  assign w_206 = w_171;
  assign w_207 = w_172;
  assign w_208 = w_173;
  assign w_209 = w_174;
  assign w_210 = w_175;
  assign w_211 = w_176;
  assign w_212 = w_177;
  assign w_213 = w_178;
  assign w_214 = w_179;
  assign w_215 = w_180;
  assign w_216 = w_181;
  assign w_217 = w_182;
  assign w_218 = w_183;
  assign w_219 = w_184;
  assign w_220 = w_185;
  assign w_221 = w_186;
  assign w_222 = w_187;
  assign w_223 = w_188;
  assign w_224 = w_189;
  assign w_225 = w_190;
  assign w_226 = w_191;
  assign w_641 = w_640;
  assign w_646 = w_645;
  assign w_651 = w_650;
  assign w_690 = w_689;
  assign w_693 = w_692;
  assign w_660 = w_657;
  assign w_661 = w_658;
  assign w_662 = w_659;
  assign w_697 = w_696;
  assign w_835 = w_834;
  assign w_843 = w_842;
  assign w_888 = w_887;
  assign w_893 = w_892;
  assign w_896 = w_895;
  assign w_883 = w_879;
  assign w_884 = w_471;
  assign w_885 = w_882;
  assign w_1324 = w_1323;
  assign w_595 = w_594;
  assign w_471 = w_457;
  assign w_472 = w_458;
  assign w_473 = w_465;
  assign w_474 = w_466;
  assign w_475 = w_467;
  assign w_476 = w_468;
  assign w_477 = w_469;
  assign w_478 = w_470;
  assign w_1362 = w_1356;
  assign w_1363 = w_1357;
  assign w_1364 = w_1358;
  assign w_1365 = w_1359;
  assign w_1366 = w_1360;
  assign w_1367 = w_1361;
  assign w_1356 = w_1343;
  assign w_1357 = w_1344;
  assign w_1358 = w_1345;
  assign w_1359 = w_1346;
  assign w_1360 = w_1347;
  assign w_1361 = w_1348;
  assign w_1369 = w_1337;
  assign w_1370 = w_1338;
  assign w_1371 = w_1339;
  assign w_1372 = w_1340;
  assign w_1373 = w_1341;
  assign w_1374 = w_1342;
  assign w_1375 = w_1362;
  assign w_1376 = w_1363;
  assign w_1377 = w_1364;
  assign w_1378 = w_1365;
  assign w_1379 = w_1366;
  assign w_1380 = w_1367;
  assign w_1337 = w_599;
  assign w_1338 = w_2;
  assign w_1339 = w_633;
  assign w_1340 = w_704;
  assign w_1341 = w_727;
  assign w_1342 = w_1297;
  assign w_1343 = w_1306;
  assign w_1344 = w_1312;
  assign w_1345 = w_1319;
  assign w_1346 = w_1321;
  assign w_1347 = w_1326;
  assign w_1348 = w_1329;
  assign w_1349 = w_1330;
  assign w_1350 = w_1331;
  assign w_1351 = w_1332;
  assign w_1352 = w_1333;
  assign w_1353 = w_1334;
  assign w_1354 = w_1335;
  assign w_465 = w_459;
  assign w_466 = w_460;
  assign w_467 = w_461;
  assign w_468 = w_462;
  assign w_469 = w_463;
  assign w_470 = w_464;
  assign w_1330 = w_459;
  assign w_1331 = w_460;
  assign w_1332 = w_461;
  assign w_1333 = w_462;
  assign w_1334 = w_463;
  assign w_1335 = w_464;
  assign w_457 = w_228;
  assign w_458 = w_423;
  assign w_1547 = w_1453;
  assign w_1548 = w_1455;
  assign w_1549 = w_1457;
  assign w_1550 = w_1459;
  assign w_1551 = w_1461;
  assign w_1552 = w_1463;
  assign w_1553 = w_1465;
  assign w_1554 = w_1467;
  assign w_1555 = w_1469;
  assign w_1556 = w_1471;
  assign w_1557 = w_1473;
  assign w_1558 = w_1475;
  assign w_1559 = w_1477;
  assign w_1560 = w_1479;
  assign w_1561 = w_1481;
  assign w_1562 = w_1483;
  assign w_1563 = w_1485;
  assign w_1564 = w_1487;
  assign w_1565 = w_1489;
  assign w_1566 = w_1491;
  assign w_1567 = w_1493;
  assign w_1568 = w_1495;
  assign w_1569 = w_1497;
  assign w_1570 = w_1499;
  assign w_1571 = w_1501;
  assign w_1572 = w_1503;
  assign w_1573 = w_1505;
  assign w_1574 = w_1507;
  assign w_1575 = w_1509;
  assign w_1576 = w_1511;
  assign w_1577 = w_1513;
  assign w_1578 = w_1451;
  assign w_1420 = w_1388;
  assign w_1421 = w_1389;
  assign w_1422 = w_1390;
  assign w_1423 = w_1391;
  assign w_1424 = w_1392;
  assign w_1425 = w_1393;
  assign w_1426 = w_1394;
  assign w_1427 = w_1395;
  assign w_1428 = w_1396;
  assign w_1429 = w_1397;
  assign w_1430 = w_1398;
  assign w_1431 = w_1399;
  assign w_1432 = w_1400;
  assign w_1433 = w_1401;
  assign w_1434 = w_1402;
  assign w_1435 = w_1403;
  assign w_1436 = w_1404;
  assign w_1437 = w_1405;
  assign w_1438 = w_1406;
  assign w_1439 = w_1407;
  assign w_1440 = w_1408;
  assign w_1441 = w_1409;
  assign w_1442 = w_1410;
  assign w_1443 = w_1411;
  assign w_1444 = w_1412;
  assign w_1445 = w_1413;
  assign w_1446 = w_1414;
  assign w_1447 = w_1415;
  assign w_1448 = w_1416;
  assign w_1449 = w_1417;
  assign w_1450 = w_1418;
  assign w_1451 = w_1419;
  assign w_1514 = w_1388;
  assign w_1515 = w_1389;
  assign w_1516 = w_1390;
  assign w_1517 = w_1391;
  assign w_1518 = w_1392;
  assign w_1519 = w_1393;
  assign w_1520 = w_1394;
  assign w_1521 = w_1395;
  assign w_1522 = w_1396;
  assign w_1523 = w_1397;
  assign w_1524 = w_1398;
  assign w_1525 = w_1399;
  assign w_1526 = w_1400;
  assign w_1527 = w_1401;
  assign w_1528 = w_1402;
  assign w_1529 = w_1403;
  assign w_1530 = w_1404;
  assign w_1531 = w_1405;
  assign w_1532 = w_1406;
  assign w_1533 = w_1407;
  assign w_1534 = w_1408;
  assign w_1535 = w_1409;
  assign w_1536 = w_1410;
  assign w_1537 = w_1411;
  assign w_1538 = w_1412;
  assign w_1539 = w_1413;
  assign w_1540 = w_1414;
  assign w_1541 = w_1415;
  assign w_1542 = w_1416;
  assign w_1543 = w_1417;
  assign w_1544 = w_1418;
  assign w_1545 = w_1419;
  assign w_1579 = w_1547;
  assign w_1580 = w_1548;
  assign w_1581 = w_1549;
  assign w_1582 = w_1550;
  assign w_1583 = w_1551;
  assign w_1584 = w_1552;
  assign w_1585 = w_1553;
  assign w_1586 = w_1554;
  assign w_1587 = w_1555;
  assign w_1588 = w_1556;
  assign w_1589 = w_1557;
  assign w_1590 = w_1558;
  assign w_1591 = w_1559;
  assign w_1592 = w_1560;
  assign w_1593 = w_1561;
  assign w_1594 = w_1562;
  assign w_1595 = w_1563;
  assign w_1596 = w_1564;
  assign w_1597 = w_1565;
  assign w_1598 = w_1566;
  assign w_1599 = w_1567;
  assign w_1600 = w_1568;
  assign w_1601 = w_1569;
  assign w_1602 = w_1570;
  assign w_1603 = w_1571;
  assign w_1604 = w_1572;
  assign w_1605 = w_1573;
  assign w_1606 = w_1574;
  assign w_1607 = w_1575;
  assign w_1608 = w_1576;
  assign w_1609 = w_1577;
  assign w_1610 = w_1578;
  assign w_1616 = w_1612;
  assign w_1617 = w_1613;
  assign w_1618 = w_1614;
  assign w_1619 = w_1615;
  assign w_1612 = w_1382;
  assign w_1613 = w_1383;
  assign w_1614 = w_1384;
  assign w_1615 = w_1385;
  assign w_1382 = w_1369;
  assign w_1383 = w_1370;
  assign w_1384 = w_1371;
  assign w_1385 = w_1372;
  assign w_1386 = w_1373;
  assign w_1387 = w_1374;
  assign w_1388 = w_424;
  assign w_1389 = w_425;
  assign w_1390 = w_426;
  assign w_1391 = w_427;
  assign w_1392 = w_428;
  assign w_1393 = w_429;
  assign w_1394 = w_430;
  assign w_1395 = w_431;
  assign w_1396 = w_432;
  assign w_1397 = w_433;
  assign w_1398 = w_434;
  assign w_1399 = w_435;
  assign w_1400 = w_436;
  assign w_1401 = w_437;
  assign w_1402 = w_438;
  assign w_1403 = w_439;
  assign w_1404 = w_440;
  assign w_1405 = w_441;
  assign w_1406 = w_442;
  assign w_1407 = w_443;
  assign w_1408 = w_444;
  assign w_1409 = w_445;
  assign w_1410 = w_446;
  assign w_1411 = w_447;
  assign w_1412 = w_448;
  assign w_1413 = w_449;
  assign w_1414 = w_450;
  assign w_1415 = w_451;
  assign w_1416 = w_452;
  assign w_1417 = w_453;
  assign w_1418 = w_454;
  assign w_1419 = w_455;
  assign w_1620 = w_1375;
  assign w_1621 = w_1376;
  assign w_1622 = w_1377;
  assign w_1623 = w_1378;
  assign w_1624 = w_1379;
  assign w_1625 = w_1380;

  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_67 (.slice_in_1(w_1), .slice_out(w_67));
  eq #(.LEN(5))
    eq_68 (.eq_in_1(w_67), .eq_in_2(5'd31), .eq_out(w_68));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_69 (.slice_in_1(w_1), .slice_out(w_69));
  eq #(.LEN(5))
    eq_70 (.eq_in_1(w_69), .eq_in_2(5'd30), .eq_out(w_70));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_71 (.slice_in_1(w_1), .slice_out(w_71));
  eq #(.LEN(5))
    eq_72 (.eq_in_1(w_71), .eq_in_2(5'd29), .eq_out(w_72));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_73 (.slice_in_1(w_1), .slice_out(w_73));
  eq #(.LEN(5))
    eq_74 (.eq_in_1(w_73), .eq_in_2(5'd28), .eq_out(w_74));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_75 (.slice_in_1(w_1), .slice_out(w_75));
  eq #(.LEN(5))
    eq_76 (.eq_in_1(w_75), .eq_in_2(5'd27), .eq_out(w_76));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_77 (.slice_in_1(w_1), .slice_out(w_77));
  eq #(.LEN(5))
    eq_78 (.eq_in_1(w_77), .eq_in_2(5'd26), .eq_out(w_78));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_79 (.slice_in_1(w_1), .slice_out(w_79));
  eq #(.LEN(5))
    eq_80 (.eq_in_1(w_79), .eq_in_2(5'd25), .eq_out(w_80));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_81 (.slice_in_1(w_1), .slice_out(w_81));
  eq #(.LEN(5))
    eq_82 (.eq_in_1(w_81), .eq_in_2(5'd24), .eq_out(w_82));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_83 (.slice_in_1(w_1), .slice_out(w_83));
  eq #(.LEN(5))
    eq_84 (.eq_in_1(w_83), .eq_in_2(5'd23), .eq_out(w_84));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_85 (.slice_in_1(w_1), .slice_out(w_85));
  eq #(.LEN(5))
    eq_86 (.eq_in_1(w_85), .eq_in_2(5'd22), .eq_out(w_86));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_87 (.slice_in_1(w_1), .slice_out(w_87));
  eq #(.LEN(5))
    eq_88 (.eq_in_1(w_87), .eq_in_2(5'd21), .eq_out(w_88));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_89 (.slice_in_1(w_1), .slice_out(w_89));
  eq #(.LEN(5))
    eq_90 (.eq_in_1(w_89), .eq_in_2(5'd20), .eq_out(w_90));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_91 (.slice_in_1(w_1), .slice_out(w_91));
  eq #(.LEN(5))
    eq_92 (.eq_in_1(w_91), .eq_in_2(5'd19), .eq_out(w_92));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_93 (.slice_in_1(w_1), .slice_out(w_93));
  eq #(.LEN(5))
    eq_94 (.eq_in_1(w_93), .eq_in_2(5'd18), .eq_out(w_94));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_95 (.slice_in_1(w_1), .slice_out(w_95));
  eq #(.LEN(5))
    eq_96 (.eq_in_1(w_95), .eq_in_2(5'd17), .eq_out(w_96));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_97 (.slice_in_1(w_1), .slice_out(w_97));
  eq #(.LEN(5))
    eq_98 (.eq_in_1(w_97), .eq_in_2(5'd16), .eq_out(w_98));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_99 (.slice_in_1(w_1), .slice_out(w_99));
  eq #(.LEN(5))
    eq_100 (.eq_in_1(w_99), .eq_in_2(5'd15), .eq_out(w_100));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_101 (.slice_in_1(w_1), .slice_out(w_101));
  eq #(.LEN(5))
    eq_102 (.eq_in_1(w_101), .eq_in_2(5'd14), .eq_out(w_102));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_103 (.slice_in_1(w_1), .slice_out(w_103));
  eq #(.LEN(5))
    eq_104 (.eq_in_1(w_103), .eq_in_2(5'd13), .eq_out(w_104));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_105 (.slice_in_1(w_1), .slice_out(w_105));
  eq #(.LEN(5))
    eq_106 (.eq_in_1(w_105), .eq_in_2(5'd12), .eq_out(w_106));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_107 (.slice_in_1(w_1), .slice_out(w_107));
  eq #(.LEN(5))
    eq_108 (.eq_in_1(w_107), .eq_in_2(5'd11), .eq_out(w_108));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_109 (.slice_in_1(w_1), .slice_out(w_109));
  eq #(.LEN(5))
    eq_110 (.eq_in_1(w_109), .eq_in_2(5'd10), .eq_out(w_110));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_111 (.slice_in_1(w_1), .slice_out(w_111));
  eq #(.LEN(5))
    eq_112 (.eq_in_1(w_111), .eq_in_2(5'd9), .eq_out(w_112));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_113 (.slice_in_1(w_1), .slice_out(w_113));
  eq #(.LEN(5))
    eq_114 (.eq_in_1(w_113), .eq_in_2(5'd8), .eq_out(w_114));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_115 (.slice_in_1(w_1), .slice_out(w_115));
  eq #(.LEN(5))
    eq_116 (.eq_in_1(w_115), .eq_in_2(5'd7), .eq_out(w_116));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_117 (.slice_in_1(w_1), .slice_out(w_117));
  eq #(.LEN(5))
    eq_118 (.eq_in_1(w_117), .eq_in_2(5'd6), .eq_out(w_118));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_119 (.slice_in_1(w_1), .slice_out(w_119));
  eq #(.LEN(5))
    eq_120 (.eq_in_1(w_119), .eq_in_2(5'd5), .eq_out(w_120));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_121 (.slice_in_1(w_1), .slice_out(w_121));
  eq #(.LEN(5))
    eq_122 (.eq_in_1(w_121), .eq_in_2(5'd4), .eq_out(w_122));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_123 (.slice_in_1(w_1), .slice_out(w_123));
  eq #(.LEN(5))
    eq_124 (.eq_in_1(w_123), .eq_in_2(5'd3), .eq_out(w_124));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_125 (.slice_in_1(w_1), .slice_out(w_125));
  eq #(.LEN(5))
    eq_126 (.eq_in_1(w_125), .eq_in_2(5'd2), .eq_out(w_126));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_127 (.slice_in_1(w_1), .slice_out(w_127));
  eq #(.LEN(5))
    eq_128 (.eq_in_1(w_127), .eq_in_2(5'd1), .eq_out(w_128));
  mux21_comp #(.LEN(32))
    mux21_comp_129 (.mux21_comp_sel(w_128), .mux21_comp_in_1(w_65), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_129));
  mux21_comp #(.LEN(32))
    mux21_comp_130 (.mux21_comp_sel(w_126), .mux21_comp_in_1(w_64), .mux21_comp_in_2(w_129), .mux21_comp_out(w_130));
  mux21_comp #(.LEN(32))
    mux21_comp_131 (.mux21_comp_sel(w_124), .mux21_comp_in_1(w_63), .mux21_comp_in_2(w_130), .mux21_comp_out(w_131));
  mux21_comp #(.LEN(32))
    mux21_comp_132 (.mux21_comp_sel(w_122), .mux21_comp_in_1(w_62), .mux21_comp_in_2(w_131), .mux21_comp_out(w_132));
  mux21_comp #(.LEN(32))
    mux21_comp_133 (.mux21_comp_sel(w_120), .mux21_comp_in_1(w_61), .mux21_comp_in_2(w_132), .mux21_comp_out(w_133));
  mux21_comp #(.LEN(32))
    mux21_comp_134 (.mux21_comp_sel(w_118), .mux21_comp_in_1(w_60), .mux21_comp_in_2(w_133), .mux21_comp_out(w_134));
  mux21_comp #(.LEN(32))
    mux21_comp_135 (.mux21_comp_sel(w_116), .mux21_comp_in_1(w_59), .mux21_comp_in_2(w_134), .mux21_comp_out(w_135));
  mux21_comp #(.LEN(32))
    mux21_comp_136 (.mux21_comp_sel(w_114), .mux21_comp_in_1(w_58), .mux21_comp_in_2(w_135), .mux21_comp_out(w_136));
  mux21_comp #(.LEN(32))
    mux21_comp_137 (.mux21_comp_sel(w_112), .mux21_comp_in_1(w_57), .mux21_comp_in_2(w_136), .mux21_comp_out(w_137));
  mux21_comp #(.LEN(32))
    mux21_comp_138 (.mux21_comp_sel(w_110), .mux21_comp_in_1(w_56), .mux21_comp_in_2(w_137), .mux21_comp_out(w_138));
  mux21_comp #(.LEN(32))
    mux21_comp_139 (.mux21_comp_sel(w_108), .mux21_comp_in_1(w_55), .mux21_comp_in_2(w_138), .mux21_comp_out(w_139));
  mux21_comp #(.LEN(32))
    mux21_comp_140 (.mux21_comp_sel(w_106), .mux21_comp_in_1(w_54), .mux21_comp_in_2(w_139), .mux21_comp_out(w_140));
  mux21_comp #(.LEN(32))
    mux21_comp_141 (.mux21_comp_sel(w_104), .mux21_comp_in_1(w_53), .mux21_comp_in_2(w_140), .mux21_comp_out(w_141));
  mux21_comp #(.LEN(32))
    mux21_comp_142 (.mux21_comp_sel(w_102), .mux21_comp_in_1(w_52), .mux21_comp_in_2(w_141), .mux21_comp_out(w_142));
  mux21_comp #(.LEN(32))
    mux21_comp_143 (.mux21_comp_sel(w_100), .mux21_comp_in_1(w_51), .mux21_comp_in_2(w_142), .mux21_comp_out(w_143));
  mux21_comp #(.LEN(32))
    mux21_comp_144 (.mux21_comp_sel(w_98), .mux21_comp_in_1(w_50), .mux21_comp_in_2(w_143), .mux21_comp_out(w_144));
  mux21_comp #(.LEN(32))
    mux21_comp_145 (.mux21_comp_sel(w_96), .mux21_comp_in_1(w_49), .mux21_comp_in_2(w_144), .mux21_comp_out(w_145));
  mux21_comp #(.LEN(32))
    mux21_comp_146 (.mux21_comp_sel(w_94), .mux21_comp_in_1(w_48), .mux21_comp_in_2(w_145), .mux21_comp_out(w_146));
  mux21_comp #(.LEN(32))
    mux21_comp_147 (.mux21_comp_sel(w_92), .mux21_comp_in_1(w_47), .mux21_comp_in_2(w_146), .mux21_comp_out(w_147));
  mux21_comp #(.LEN(32))
    mux21_comp_148 (.mux21_comp_sel(w_90), .mux21_comp_in_1(w_46), .mux21_comp_in_2(w_147), .mux21_comp_out(w_148));
  mux21_comp #(.LEN(32))
    mux21_comp_149 (.mux21_comp_sel(w_88), .mux21_comp_in_1(w_45), .mux21_comp_in_2(w_148), .mux21_comp_out(w_149));
  mux21_comp #(.LEN(32))
    mux21_comp_150 (.mux21_comp_sel(w_86), .mux21_comp_in_1(w_44), .mux21_comp_in_2(w_149), .mux21_comp_out(w_150));
  mux21_comp #(.LEN(32))
    mux21_comp_151 (.mux21_comp_sel(w_84), .mux21_comp_in_1(w_43), .mux21_comp_in_2(w_150), .mux21_comp_out(w_151));
  mux21_comp #(.LEN(32))
    mux21_comp_152 (.mux21_comp_sel(w_82), .mux21_comp_in_1(w_42), .mux21_comp_in_2(w_151), .mux21_comp_out(w_152));
  mux21_comp #(.LEN(32))
    mux21_comp_153 (.mux21_comp_sel(w_80), .mux21_comp_in_1(w_41), .mux21_comp_in_2(w_152), .mux21_comp_out(w_153));
  mux21_comp #(.LEN(32))
    mux21_comp_154 (.mux21_comp_sel(w_78), .mux21_comp_in_1(w_40), .mux21_comp_in_2(w_153), .mux21_comp_out(w_154));
  mux21_comp #(.LEN(32))
    mux21_comp_155 (.mux21_comp_sel(w_76), .mux21_comp_in_1(w_39), .mux21_comp_in_2(w_154), .mux21_comp_out(w_155));
  mux21_comp #(.LEN(32))
    mux21_comp_156 (.mux21_comp_sel(w_74), .mux21_comp_in_1(w_38), .mux21_comp_in_2(w_155), .mux21_comp_out(w_156));
  mux21_comp #(.LEN(32))
    mux21_comp_157 (.mux21_comp_sel(w_72), .mux21_comp_in_1(w_37), .mux21_comp_in_2(w_156), .mux21_comp_out(w_157));
  mux21_comp #(.LEN(32))
    mux21_comp_158 (.mux21_comp_sel(w_70), .mux21_comp_in_1(w_36), .mux21_comp_in_2(w_157), .mux21_comp_out(w_158));
  mux21_comp #(.LEN(32))
    mux21_comp_159 (.mux21_comp_sel(w_68), .mux21_comp_in_1(w_35), .mux21_comp_in_2(w_158), .mux21_comp_out(w_159));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_194 (.slice_in_1(w_1), .slice_out(w_194));
  eq #(.LEN(5))
    eq_328 (.eq_in_1(w_263), .eq_in_2(5'd31), .eq_out(w_328));
  eq #(.LEN(5))
    eq_329 (.eq_in_1(w_263), .eq_in_2(5'd30), .eq_out(w_329));
  eq #(.LEN(5))
    eq_330 (.eq_in_1(w_263), .eq_in_2(5'd29), .eq_out(w_330));
  eq #(.LEN(5))
    eq_331 (.eq_in_1(w_263), .eq_in_2(5'd28), .eq_out(w_331));
  eq #(.LEN(5))
    eq_332 (.eq_in_1(w_263), .eq_in_2(5'd27), .eq_out(w_332));
  eq #(.LEN(5))
    eq_333 (.eq_in_1(w_263), .eq_in_2(5'd26), .eq_out(w_333));
  eq #(.LEN(5))
    eq_334 (.eq_in_1(w_263), .eq_in_2(5'd25), .eq_out(w_334));
  eq #(.LEN(5))
    eq_335 (.eq_in_1(w_263), .eq_in_2(5'd24), .eq_out(w_335));
  eq #(.LEN(5))
    eq_336 (.eq_in_1(w_263), .eq_in_2(5'd23), .eq_out(w_336));
  eq #(.LEN(5))
    eq_337 (.eq_in_1(w_263), .eq_in_2(5'd22), .eq_out(w_337));
  eq #(.LEN(5))
    eq_338 (.eq_in_1(w_263), .eq_in_2(5'd21), .eq_out(w_338));
  eq #(.LEN(5))
    eq_339 (.eq_in_1(w_263), .eq_in_2(5'd20), .eq_out(w_339));
  eq #(.LEN(5))
    eq_340 (.eq_in_1(w_263), .eq_in_2(5'd19), .eq_out(w_340));
  eq #(.LEN(5))
    eq_341 (.eq_in_1(w_263), .eq_in_2(5'd18), .eq_out(w_341));
  eq #(.LEN(5))
    eq_342 (.eq_in_1(w_263), .eq_in_2(5'd17), .eq_out(w_342));
  eq #(.LEN(5))
    eq_343 (.eq_in_1(w_263), .eq_in_2(5'd16), .eq_out(w_343));
  eq #(.LEN(5))
    eq_344 (.eq_in_1(w_263), .eq_in_2(5'd15), .eq_out(w_344));
  eq #(.LEN(5))
    eq_345 (.eq_in_1(w_263), .eq_in_2(5'd14), .eq_out(w_345));
  eq #(.LEN(5))
    eq_346 (.eq_in_1(w_263), .eq_in_2(5'd13), .eq_out(w_346));
  eq #(.LEN(5))
    eq_347 (.eq_in_1(w_263), .eq_in_2(5'd12), .eq_out(w_347));
  eq #(.LEN(5))
    eq_348 (.eq_in_1(w_263), .eq_in_2(5'd11), .eq_out(w_348));
  eq #(.LEN(5))
    eq_349 (.eq_in_1(w_263), .eq_in_2(5'd10), .eq_out(w_349));
  eq #(.LEN(5))
    eq_350 (.eq_in_1(w_263), .eq_in_2(5'd9), .eq_out(w_350));
  eq #(.LEN(5))
    eq_351 (.eq_in_1(w_263), .eq_in_2(5'd8), .eq_out(w_351));
  eq #(.LEN(5))
    eq_352 (.eq_in_1(w_263), .eq_in_2(5'd7), .eq_out(w_352));
  eq #(.LEN(5))
    eq_353 (.eq_in_1(w_263), .eq_in_2(5'd6), .eq_out(w_353));
  eq #(.LEN(5))
    eq_354 (.eq_in_1(w_263), .eq_in_2(5'd5), .eq_out(w_354));
  eq #(.LEN(5))
    eq_355 (.eq_in_1(w_263), .eq_in_2(5'd4), .eq_out(w_355));
  eq #(.LEN(5))
    eq_356 (.eq_in_1(w_263), .eq_in_2(5'd3), .eq_out(w_356));
  eq #(.LEN(5))
    eq_357 (.eq_in_1(w_263), .eq_in_2(5'd2), .eq_out(w_357));
  eq #(.LEN(5))
    eq_358 (.eq_in_1(w_263), .eq_in_2(5'd1), .eq_out(w_358));
  mux21_comp #(.LEN(32))
    mux21_comp_359 (.mux21_comp_sel(w_358), .mux21_comp_in_1(w_326), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_359));
  mux21_comp #(.LEN(32))
    mux21_comp_360 (.mux21_comp_sel(w_357), .mux21_comp_in_1(w_325), .mux21_comp_in_2(w_359), .mux21_comp_out(w_360));
  mux21_comp #(.LEN(32))
    mux21_comp_361 (.mux21_comp_sel(w_356), .mux21_comp_in_1(w_324), .mux21_comp_in_2(w_360), .mux21_comp_out(w_361));
  mux21_comp #(.LEN(32))
    mux21_comp_362 (.mux21_comp_sel(w_355), .mux21_comp_in_1(w_323), .mux21_comp_in_2(w_361), .mux21_comp_out(w_362));
  mux21_comp #(.LEN(32))
    mux21_comp_363 (.mux21_comp_sel(w_354), .mux21_comp_in_1(w_322), .mux21_comp_in_2(w_362), .mux21_comp_out(w_363));
  mux21_comp #(.LEN(32))
    mux21_comp_364 (.mux21_comp_sel(w_353), .mux21_comp_in_1(w_321), .mux21_comp_in_2(w_363), .mux21_comp_out(w_364));
  mux21_comp #(.LEN(32))
    mux21_comp_365 (.mux21_comp_sel(w_352), .mux21_comp_in_1(w_320), .mux21_comp_in_2(w_364), .mux21_comp_out(w_365));
  mux21_comp #(.LEN(32))
    mux21_comp_366 (.mux21_comp_sel(w_351), .mux21_comp_in_1(w_319), .mux21_comp_in_2(w_365), .mux21_comp_out(w_366));
  mux21_comp #(.LEN(32))
    mux21_comp_367 (.mux21_comp_sel(w_350), .mux21_comp_in_1(w_318), .mux21_comp_in_2(w_366), .mux21_comp_out(w_367));
  mux21_comp #(.LEN(32))
    mux21_comp_368 (.mux21_comp_sel(w_349), .mux21_comp_in_1(w_317), .mux21_comp_in_2(w_367), .mux21_comp_out(w_368));
  mux21_comp #(.LEN(32))
    mux21_comp_369 (.mux21_comp_sel(w_348), .mux21_comp_in_1(w_316), .mux21_comp_in_2(w_368), .mux21_comp_out(w_369));
  mux21_comp #(.LEN(32))
    mux21_comp_370 (.mux21_comp_sel(w_347), .mux21_comp_in_1(w_315), .mux21_comp_in_2(w_369), .mux21_comp_out(w_370));
  mux21_comp #(.LEN(32))
    mux21_comp_371 (.mux21_comp_sel(w_346), .mux21_comp_in_1(w_314), .mux21_comp_in_2(w_370), .mux21_comp_out(w_371));
  mux21_comp #(.LEN(32))
    mux21_comp_372 (.mux21_comp_sel(w_345), .mux21_comp_in_1(w_313), .mux21_comp_in_2(w_371), .mux21_comp_out(w_372));
  mux21_comp #(.LEN(32))
    mux21_comp_373 (.mux21_comp_sel(w_344), .mux21_comp_in_1(w_312), .mux21_comp_in_2(w_372), .mux21_comp_out(w_373));
  mux21_comp #(.LEN(32))
    mux21_comp_374 (.mux21_comp_sel(w_343), .mux21_comp_in_1(w_311), .mux21_comp_in_2(w_373), .mux21_comp_out(w_374));
  mux21_comp #(.LEN(32))
    mux21_comp_375 (.mux21_comp_sel(w_342), .mux21_comp_in_1(w_310), .mux21_comp_in_2(w_374), .mux21_comp_out(w_375));
  mux21_comp #(.LEN(32))
    mux21_comp_376 (.mux21_comp_sel(w_341), .mux21_comp_in_1(w_309), .mux21_comp_in_2(w_375), .mux21_comp_out(w_376));
  mux21_comp #(.LEN(32))
    mux21_comp_377 (.mux21_comp_sel(w_340), .mux21_comp_in_1(w_308), .mux21_comp_in_2(w_376), .mux21_comp_out(w_377));
  mux21_comp #(.LEN(32))
    mux21_comp_378 (.mux21_comp_sel(w_339), .mux21_comp_in_1(w_307), .mux21_comp_in_2(w_377), .mux21_comp_out(w_378));
  mux21_comp #(.LEN(32))
    mux21_comp_379 (.mux21_comp_sel(w_338), .mux21_comp_in_1(w_306), .mux21_comp_in_2(w_378), .mux21_comp_out(w_379));
  mux21_comp #(.LEN(32))
    mux21_comp_380 (.mux21_comp_sel(w_337), .mux21_comp_in_1(w_305), .mux21_comp_in_2(w_379), .mux21_comp_out(w_380));
  mux21_comp #(.LEN(32))
    mux21_comp_381 (.mux21_comp_sel(w_336), .mux21_comp_in_1(w_304), .mux21_comp_in_2(w_380), .mux21_comp_out(w_381));
  mux21_comp #(.LEN(32))
    mux21_comp_382 (.mux21_comp_sel(w_335), .mux21_comp_in_1(w_303), .mux21_comp_in_2(w_381), .mux21_comp_out(w_382));
  mux21_comp #(.LEN(32))
    mux21_comp_383 (.mux21_comp_sel(w_334), .mux21_comp_in_1(w_302), .mux21_comp_in_2(w_382), .mux21_comp_out(w_383));
  mux21_comp #(.LEN(32))
    mux21_comp_384 (.mux21_comp_sel(w_333), .mux21_comp_in_1(w_301), .mux21_comp_in_2(w_383), .mux21_comp_out(w_384));
  mux21_comp #(.LEN(32))
    mux21_comp_385 (.mux21_comp_sel(w_332), .mux21_comp_in_1(w_300), .mux21_comp_in_2(w_384), .mux21_comp_out(w_385));
  mux21_comp #(.LEN(32))
    mux21_comp_386 (.mux21_comp_sel(w_331), .mux21_comp_in_1(w_299), .mux21_comp_in_2(w_385), .mux21_comp_out(w_386));
  mux21_comp #(.LEN(32))
    mux21_comp_387 (.mux21_comp_sel(w_330), .mux21_comp_in_1(w_298), .mux21_comp_in_2(w_386), .mux21_comp_out(w_387));
  mux21_comp #(.LEN(32))
    mux21_comp_388 (.mux21_comp_sel(w_329), .mux21_comp_in_1(w_297), .mux21_comp_in_2(w_387), .mux21_comp_out(w_388));
  mux21_comp #(.LEN(32))
    mux21_comp_389 (.mux21_comp_sel(w_328), .mux21_comp_in_1(w_296), .mux21_comp_in_2(w_388), .mux21_comp_out(w_389));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_479 (.slice_in_1(w_1), .slice_out(w_479));
  eq #(.LEN(7))
    eq_480 (.eq_in_1(w_479), .eq_in_2(7'd19), .eq_out(w_480));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_481 (.slice_in_1(w_1), .slice_out(w_481));
  eq #(.LEN(7))
    eq_482 (.eq_in_1(w_481), .eq_in_2(7'd3), .eq_out(w_482));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_483 (.slice_in_1(w_1), .slice_out(w_483));
  eq #(.LEN(7))
    eq_484 (.eq_in_1(w_483), .eq_in_2(7'd103), .eq_out(w_484));
  or_comp #(.LEN(1))
    or_comp_485 (.or_comp_in_1(w_482), .or_comp_in_2(w_484), .or_comp_out(w_485));
  or_comp #(.LEN(1))
    or_comp_486 (.or_comp_in_1(w_480), .or_comp_in_2(w_485), .or_comp_out(w_486));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_487 (.slice_in_1(w_1), .slice_out(w_487));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_488 (.slice_in_1(w_1), .slice_out(w_488));
  concat #(.LEN1(7), .LEN2(5))
    concat_489 (.concat_in_1(w_487), .concat_in_2(w_488), .concat_out(w_489));
  slice #(.LEN(12), .LOWER(11), .UPPER(12))
    slice_490 (.slice_in_1(w_489), .slice_out(w_490));
  not_comp #(.LEN(20))
    not_comp_491 (.not_comp_in_1(20'd0), .not_comp_out(w_491));
  mux21_comp #(.LEN(20))
    mux21_comp_492 (.mux21_comp_sel(w_490), .mux21_comp_in_1(w_491), .mux21_comp_in_2(20'd0), .mux21_comp_out(w_492));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_493 (.slice_in_1(w_1), .slice_out(w_493));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_494 (.slice_in_1(w_1), .slice_out(w_494));
  concat #(.LEN1(7), .LEN2(5))
    concat_495 (.concat_in_1(w_493), .concat_in_2(w_494), .concat_out(w_495));
  concat #(.LEN1(20), .LEN2(12))
    concat_496 (.concat_in_1(w_492), .concat_in_2(w_495), .concat_out(w_496));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_497 (.slice_in_1(w_1), .slice_out(w_497));
  eq #(.LEN(7))
    eq_498 (.eq_in_1(w_497), .eq_in_2(7'd35), .eq_out(w_498));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_499 (.slice_in_1(w_1), .slice_out(w_499));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_500 (.slice_in_1(w_1), .slice_out(w_500));
  concat #(.LEN1(7), .LEN2(5))
    concat_501 (.concat_in_1(w_499), .concat_in_2(w_500), .concat_out(w_501));
  slice #(.LEN(12), .LOWER(11), .UPPER(12))
    slice_502 (.slice_in_1(w_501), .slice_out(w_502));
  not_comp #(.LEN(20))
    not_comp_503 (.not_comp_in_1(20'd0), .not_comp_out(w_503));
  mux21_comp #(.LEN(20))
    mux21_comp_504 (.mux21_comp_sel(w_502), .mux21_comp_in_1(w_503), .mux21_comp_in_2(20'd0), .mux21_comp_out(w_504));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_505 (.slice_in_1(w_1), .slice_out(w_505));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_506 (.slice_in_1(w_1), .slice_out(w_506));
  concat #(.LEN1(7), .LEN2(5))
    concat_507 (.concat_in_1(w_505), .concat_in_2(w_506), .concat_out(w_507));
  concat #(.LEN1(20), .LEN2(12))
    concat_508 (.concat_in_1(w_504), .concat_in_2(w_507), .concat_out(w_508));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_509 (.slice_in_1(w_1), .slice_out(w_509));
  eq #(.LEN(7))
    eq_510 (.eq_in_1(w_509), .eq_in_2(7'd99), .eq_out(w_510));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_511 (.slice_in_1(w_1), .slice_out(w_511));
  slice #(.LEN(7), .LOWER(6), .UPPER(7))
    slice_512 (.slice_in_1(w_511), .slice_out(w_512));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_513 (.slice_in_1(w_1), .slice_out(w_513));
  slice #(.LEN(5), .LOWER(0), .UPPER(1))
    slice_514 (.slice_in_1(w_513), .slice_out(w_514));
  concat #(.LEN1(1), .LEN2(1))
    concat_515 (.concat_in_1(w_512), .concat_in_2(w_514), .concat_out(w_515));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_516 (.slice_in_1(w_1), .slice_out(w_516));
  slice #(.LEN(7), .LOWER(0), .UPPER(6))
    slice_517 (.slice_in_1(w_516), .slice_out(w_517));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_518 (.slice_in_1(w_1), .slice_out(w_518));
  not_comp #(.LEN(5))
    not_comp_519 (.not_comp_in_1(5'd1), .not_comp_out(w_519));
  and_comp #(.LEN(5))
    and_comp_520 (.and_comp_in_1(w_518), .and_comp_in_2(w_519), .and_comp_out(w_520));
  concat #(.LEN1(6), .LEN2(5))
    concat_521 (.concat_in_1(w_517), .concat_in_2(w_520), .concat_out(w_521));
  concat #(.LEN1(2), .LEN2(11))
    concat_522 (.concat_in_1(w_515), .concat_in_2(w_521), .concat_out(w_522));
  slice #(.LEN(13), .LOWER(12), .UPPER(13))
    slice_523 (.slice_in_1(w_522), .slice_out(w_523));
  not_comp #(.LEN(19))
    not_comp_524 (.not_comp_in_1(19'd0), .not_comp_out(w_524));
  mux21_comp #(.LEN(19))
    mux21_comp_525 (.mux21_comp_sel(w_523), .mux21_comp_in_1(w_524), .mux21_comp_in_2(19'd0), .mux21_comp_out(w_525));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_526 (.slice_in_1(w_1), .slice_out(w_526));
  slice #(.LEN(7), .LOWER(6), .UPPER(7))
    slice_527 (.slice_in_1(w_526), .slice_out(w_527));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_528 (.slice_in_1(w_1), .slice_out(w_528));
  slice #(.LEN(5), .LOWER(0), .UPPER(1))
    slice_529 (.slice_in_1(w_528), .slice_out(w_529));
  concat #(.LEN1(1), .LEN2(1))
    concat_530 (.concat_in_1(w_527), .concat_in_2(w_529), .concat_out(w_530));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_531 (.slice_in_1(w_1), .slice_out(w_531));
  slice #(.LEN(7), .LOWER(0), .UPPER(6))
    slice_532 (.slice_in_1(w_531), .slice_out(w_532));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_533 (.slice_in_1(w_1), .slice_out(w_533));
  not_comp #(.LEN(5))
    not_comp_534 (.not_comp_in_1(5'd1), .not_comp_out(w_534));
  and_comp #(.LEN(5))
    and_comp_535 (.and_comp_in_1(w_533), .and_comp_in_2(w_534), .and_comp_out(w_535));
  concat #(.LEN1(6), .LEN2(5))
    concat_536 (.concat_in_1(w_532), .concat_in_2(w_535), .concat_out(w_536));
  concat #(.LEN1(2), .LEN2(11))
    concat_537 (.concat_in_1(w_530), .concat_in_2(w_536), .concat_out(w_537));
  concat #(.LEN1(19), .LEN2(13))
    concat_538 (.concat_in_1(w_525), .concat_in_2(w_537), .concat_out(w_538));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_539 (.slice_in_1(w_1), .slice_out(w_539));
  eq #(.LEN(7))
    eq_540 (.eq_in_1(w_539), .eq_in_2(7'd55), .eq_out(w_540));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_541 (.slice_in_1(w_1), .slice_out(w_541));
  eq #(.LEN(7))
    eq_542 (.eq_in_1(w_541), .eq_in_2(7'd23), .eq_out(w_542));
  or_comp #(.LEN(1))
    or_comp_543 (.or_comp_in_1(w_540), .or_comp_in_2(w_542), .or_comp_out(w_543));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_544 (.slice_in_1(w_1), .slice_out(w_544));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_545 (.slice_in_1(w_1), .slice_out(w_545));
  concat #(.LEN1(7), .LEN2(5))
    concat_546 (.concat_in_1(w_544), .concat_in_2(w_545), .concat_out(w_546));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_547 (.slice_in_1(w_1), .slice_out(w_547));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_548 (.slice_in_1(w_1), .slice_out(w_548));
  concat #(.LEN1(5), .LEN2(3))
    concat_549 (.concat_in_1(w_547), .concat_in_2(w_548), .concat_out(w_549));
  concat #(.LEN1(12), .LEN2(8))
    concat_550 (.concat_in_1(w_546), .concat_in_2(w_549), .concat_out(w_550));
  concat #(.LEN1(20), .LEN2(12))
    concat_551 (.concat_in_1(w_550), .concat_in_2(12'd0), .concat_out(w_551));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_552 (.slice_in_1(w_1), .slice_out(w_552));
  eq #(.LEN(7))
    eq_553 (.eq_in_1(w_552), .eq_in_2(7'd111), .eq_out(w_553));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_554 (.slice_in_1(w_1), .slice_out(w_554));
  slice #(.LEN(7), .LOWER(6), .UPPER(7))
    slice_555 (.slice_in_1(w_554), .slice_out(w_555));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_556 (.slice_in_1(w_1), .slice_out(w_556));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_557 (.slice_in_1(w_1), .slice_out(w_557));
  concat #(.LEN1(5), .LEN2(3))
    concat_558 (.concat_in_1(w_556), .concat_in_2(w_557), .concat_out(w_558));
  concat #(.LEN1(1), .LEN2(8))
    concat_559 (.concat_in_1(w_555), .concat_in_2(w_558), .concat_out(w_559));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_560 (.slice_in_1(w_1), .slice_out(w_560));
  slice #(.LEN(5), .LOWER(0), .UPPER(1))
    slice_561 (.slice_in_1(w_560), .slice_out(w_561));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_562 (.slice_in_1(w_1), .slice_out(w_562));
  slice #(.LEN(7), .LOWER(0), .UPPER(6))
    slice_563 (.slice_in_1(w_562), .slice_out(w_563));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_564 (.slice_in_1(w_1), .slice_out(w_564));
  not_comp #(.LEN(5))
    not_comp_565 (.not_comp_in_1(5'd1), .not_comp_out(w_565));
  and_comp #(.LEN(5))
    and_comp_566 (.and_comp_in_1(w_564), .and_comp_in_2(w_565), .and_comp_out(w_566));
  concat #(.LEN1(6), .LEN2(5))
    concat_567 (.concat_in_1(w_563), .concat_in_2(w_566), .concat_out(w_567));
  concat #(.LEN1(1), .LEN2(11))
    concat_568 (.concat_in_1(w_561), .concat_in_2(w_567), .concat_out(w_568));
  concat #(.LEN1(9), .LEN2(12))
    concat_569 (.concat_in_1(w_559), .concat_in_2(w_568), .concat_out(w_569));
  slice #(.LEN(21), .LOWER(20), .UPPER(21))
    slice_570 (.slice_in_1(w_569), .slice_out(w_570));
  not_comp #(.LEN(11))
    not_comp_571 (.not_comp_in_1(11'd0), .not_comp_out(w_571));
  mux21_comp #(.LEN(11))
    mux21_comp_572 (.mux21_comp_sel(w_570), .mux21_comp_in_1(w_571), .mux21_comp_in_2(11'd0), .mux21_comp_out(w_572));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_573 (.slice_in_1(w_1), .slice_out(w_573));
  slice #(.LEN(7), .LOWER(6), .UPPER(7))
    slice_574 (.slice_in_1(w_573), .slice_out(w_574));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_575 (.slice_in_1(w_1), .slice_out(w_575));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_576 (.slice_in_1(w_1), .slice_out(w_576));
  concat #(.LEN1(5), .LEN2(3))
    concat_577 (.concat_in_1(w_575), .concat_in_2(w_576), .concat_out(w_577));
  concat #(.LEN1(1), .LEN2(8))
    concat_578 (.concat_in_1(w_574), .concat_in_2(w_577), .concat_out(w_578));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_579 (.slice_in_1(w_1), .slice_out(w_579));
  slice #(.LEN(5), .LOWER(0), .UPPER(1))
    slice_580 (.slice_in_1(w_579), .slice_out(w_580));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_581 (.slice_in_1(w_1), .slice_out(w_581));
  slice #(.LEN(7), .LOWER(0), .UPPER(6))
    slice_582 (.slice_in_1(w_581), .slice_out(w_582));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_583 (.slice_in_1(w_1), .slice_out(w_583));
  not_comp #(.LEN(5))
    not_comp_584 (.not_comp_in_1(5'd1), .not_comp_out(w_584));
  and_comp #(.LEN(5))
    and_comp_585 (.and_comp_in_1(w_583), .and_comp_in_2(w_584), .and_comp_out(w_585));
  concat #(.LEN1(6), .LEN2(5))
    concat_586 (.concat_in_1(w_582), .concat_in_2(w_585), .concat_out(w_586));
  concat #(.LEN1(1), .LEN2(11))
    concat_587 (.concat_in_1(w_580), .concat_in_2(w_586), .concat_out(w_587));
  concat #(.LEN1(9), .LEN2(12))
    concat_588 (.concat_in_1(w_578), .concat_in_2(w_587), .concat_out(w_588));
  concat #(.LEN1(11), .LEN2(21))
    concat_589 (.concat_in_1(w_572), .concat_in_2(w_588), .concat_out(w_589));
  mux21_comp #(.LEN(32))
    mux21_comp_590 (.mux21_comp_sel(w_553), .mux21_comp_in_1(w_589), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_590));
  mux21_comp #(.LEN(32))
    mux21_comp_591 (.mux21_comp_sel(w_543), .mux21_comp_in_1(w_551), .mux21_comp_in_2(w_590), .mux21_comp_out(w_591));
  mux21_comp #(.LEN(32))
    mux21_comp_592 (.mux21_comp_sel(w_510), .mux21_comp_in_1(w_538), .mux21_comp_in_2(w_591), .mux21_comp_out(w_592));
  mux21_comp #(.LEN(32))
    mux21_comp_593 (.mux21_comp_sel(w_498), .mux21_comp_in_1(w_508), .mux21_comp_in_2(w_592), .mux21_comp_out(w_593));
  mux21_comp #(.LEN(32))
    mux21_comp_594 (.mux21_comp_sel(w_486), .mux21_comp_in_1(w_496), .mux21_comp_in_2(w_593), .mux21_comp_out(w_594));
  not_comp #(.LEN(1))
    not_comp_596 (.not_comp_in_1(w_0), .not_comp_out(w_596));
  mux21_comp #(.LEN(1))
    mux21_comp_597 (.mux21_comp_sel(w_474), .mux21_comp_in_1(1'd1), .mux21_comp_in_2(1'd0), .mux21_comp_out(w_597));
  mux21_comp #(.LEN(1))
    mux21_comp_598 (.mux21_comp_sel(w_473), .mux21_comp_in_1(w_597), .mux21_comp_in_2(1'd0), .mux21_comp_out(w_598));
  mux21_comp #(.LEN(1))
    mux21_comp_599 (.mux21_comp_sel(w_596), .mux21_comp_in_1(1'd0), .mux21_comp_in_2(w_598), .mux21_comp_out(w_599));
  eq #(.LEN(3))
    eq_600 (.eq_in_1(w_478), .eq_in_2(3'd1), .eq_out(w_600));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_601 (.slice_in_1(w_1), .slice_out(w_601));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_602 (.slice_in_1(w_1), .slice_out(w_602));
  concat #(.LEN1(7), .LEN2(5))
    concat_603 (.concat_in_1(w_601), .concat_in_2(w_602), .concat_out(w_603));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_604 (.slice_in_1(w_1), .slice_out(w_604));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_605 (.slice_in_1(w_1), .slice_out(w_605));
  concat #(.LEN1(5), .LEN2(3))
    concat_606 (.concat_in_1(w_604), .concat_in_2(w_605), .concat_out(w_606));
  concat #(.LEN1(12), .LEN2(8))
    concat_607 (.concat_in_1(w_603), .concat_in_2(w_606), .concat_out(w_607));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_608 (.slice_in_1(w_1), .slice_out(w_608));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_609 (.slice_in_1(w_1), .slice_out(w_609));
  concat #(.LEN1(5), .LEN2(7))
    concat_610 (.concat_in_1(w_608), .concat_in_2(w_609), .concat_out(w_610));
  concat #(.LEN1(20), .LEN2(12))
    concat_611 (.concat_in_1(w_607), .concat_in_2(w_610), .concat_out(w_611));
  slice #(.LEN(32), .LOWER(16), .UPPER(32))
    slice_612 (.slice_in_1(w_611), .slice_out(w_612));
  slice #(.LEN(32), .LOWER(0), .UPPER(16))
    slice_613 (.slice_in_1(w_476), .slice_out(w_613));
  concat #(.LEN1(16), .LEN2(16))
    concat_614 (.concat_in_1(w_612), .concat_in_2(w_613), .concat_out(w_614));
  eq #(.LEN(3))
    eq_615 (.eq_in_1(w_478), .eq_in_2(3'd0), .eq_out(w_615));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_616 (.slice_in_1(w_1), .slice_out(w_616));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_617 (.slice_in_1(w_1), .slice_out(w_617));
  concat #(.LEN1(7), .LEN2(5))
    concat_618 (.concat_in_1(w_616), .concat_in_2(w_617), .concat_out(w_618));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_619 (.slice_in_1(w_1), .slice_out(w_619));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_620 (.slice_in_1(w_1), .slice_out(w_620));
  concat #(.LEN1(5), .LEN2(3))
    concat_621 (.concat_in_1(w_619), .concat_in_2(w_620), .concat_out(w_621));
  concat #(.LEN1(12), .LEN2(8))
    concat_622 (.concat_in_1(w_618), .concat_in_2(w_621), .concat_out(w_622));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_623 (.slice_in_1(w_1), .slice_out(w_623));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_624 (.slice_in_1(w_1), .slice_out(w_624));
  concat #(.LEN1(5), .LEN2(7))
    concat_625 (.concat_in_1(w_623), .concat_in_2(w_624), .concat_out(w_625));
  concat #(.LEN1(20), .LEN2(12))
    concat_626 (.concat_in_1(w_622), .concat_in_2(w_625), .concat_out(w_626));
  slice #(.LEN(32), .LOWER(8), .UPPER(32))
    slice_627 (.slice_in_1(w_626), .slice_out(w_627));
  slice #(.LEN(32), .LOWER(0), .UPPER(8))
    slice_628 (.slice_in_1(w_476), .slice_out(w_628));
  concat #(.LEN1(24), .LEN2(8))
    concat_629 (.concat_in_1(w_627), .concat_in_2(w_628), .concat_out(w_629));
  mux21_comp #(.LEN(32))
    mux21_comp_630 (.mux21_comp_sel(w_615), .mux21_comp_in_1(w_629), .mux21_comp_in_2(w_476), .mux21_comp_out(w_630));
  mux21_comp #(.LEN(32))
    mux21_comp_631 (.mux21_comp_sel(w_600), .mux21_comp_in_1(w_614), .mux21_comp_in_2(w_630), .mux21_comp_out(w_631));
  mux21_comp #(.LEN(32))
    mux21_comp_632 (.mux21_comp_sel(w_474), .mux21_comp_in_1(w_631), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_632));
  mux21_comp #(.LEN(32))
    mux21_comp_633 (.mux21_comp_sel(w_473), .mux21_comp_in_1(w_632), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_633));
  not_comp #(.LEN(1))
    not_comp_634 (.not_comp_in_1(w_0), .not_comp_out(w_634));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_635 (.slice_in_1(w_1), .slice_out(w_635));
  eq #(.LEN(7))
    eq_636 (.eq_in_1(w_635), .eq_in_2(7'd35), .eq_out(w_636));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_637 (.slice_in_1(w_1), .slice_out(w_637));
  eq #(.LEN(7))
    eq_638 (.eq_in_1(w_637), .eq_in_2(7'd3), .eq_out(w_638));
  or_comp #(.LEN(1))
    or_comp_639 (.or_comp_in_1(w_636), .or_comp_in_2(w_638), .or_comp_out(w_639));
  add #(.LEN(32))
    add_640 (.add_in_1(w_471), .add_in_2(w_595), .add_out(w_640));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_642 (.slice_in_1(w_641), .slice_out(w_642));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_643 (.slice_in_1(w_1), .slice_out(w_643));
  eq #(.LEN(7))
    eq_644 (.eq_in_1(w_643), .eq_in_2(7'd111), .eq_out(w_644));
  add #(.LEN(32))
    add_645 (.add_in_1(w_2), .add_in_2(w_595), .add_out(w_645));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_647 (.slice_in_1(w_646), .slice_out(w_647));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_648 (.slice_in_1(w_1), .slice_out(w_648));
  eq #(.LEN(7))
    eq_649 (.eq_in_1(w_648), .eq_in_2(7'd103), .eq_out(w_649));
  add #(.LEN(32))
    add_650 (.add_in_1(w_471), .add_in_2(w_595), .add_out(w_650));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_652 (.slice_in_1(w_651), .slice_out(w_652));
  not_comp #(.LEN(32))
    not_comp_653 (.not_comp_in_1(32'd1), .not_comp_out(w_653));
  and_comp #(.LEN(32))
    and_comp_654 (.and_comp_in_1(w_652), .and_comp_in_2(w_653), .and_comp_out(w_654));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_655 (.slice_in_1(w_1), .slice_out(w_655));
  eq #(.LEN(7))
    eq_656 (.eq_in_1(w_655), .eq_in_2(7'd99), .eq_out(w_656));
  eq #(.LEN(32))
    eq_657 (.eq_in_1(w_471), .eq_in_2(w_472), .eq_out(w_657));
  lt #(.LEN(32))
    lt_658 (.lt_in_1(w_471), .lt_in_2(w_472), .lt_out(w_658));
  ltu #(.LEN(32))
    ltu_659 (.ltu_in_1(w_471), .ltu_in_2(w_472), .ltu_out(w_659));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_663 (.slice_in_1(w_1), .slice_out(w_663));
  eq #(.LEN(3))
    eq_664 (.eq_in_1(w_663), .eq_in_2(3'd0), .eq_out(w_664));
  and_comp #(.LEN(1))
    and_comp_665 (.and_comp_in_1(w_664), .and_comp_in_2(w_660), .and_comp_out(w_665));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_666 (.slice_in_1(w_1), .slice_out(w_666));
  eq #(.LEN(3))
    eq_667 (.eq_in_1(w_666), .eq_in_2(3'd1), .eq_out(w_667));
  not_comp #(.LEN(1))
    not_comp_668 (.not_comp_in_1(w_660), .not_comp_out(w_668));
  and_comp #(.LEN(1))
    and_comp_669 (.and_comp_in_1(w_667), .and_comp_in_2(w_668), .and_comp_out(w_669));
  or_comp #(.LEN(1))
    or_comp_670 (.or_comp_in_1(w_665), .or_comp_in_2(w_669), .or_comp_out(w_670));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_671 (.slice_in_1(w_1), .slice_out(w_671));
  eq #(.LEN(3))
    eq_672 (.eq_in_1(w_671), .eq_in_2(3'd4), .eq_out(w_672));
  and_comp #(.LEN(1))
    and_comp_673 (.and_comp_in_1(w_672), .and_comp_in_2(w_661), .and_comp_out(w_673));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_674 (.slice_in_1(w_1), .slice_out(w_674));
  eq #(.LEN(3))
    eq_675 (.eq_in_1(w_674), .eq_in_2(3'd5), .eq_out(w_675));
  not_comp #(.LEN(1))
    not_comp_676 (.not_comp_in_1(w_661), .not_comp_out(w_676));
  and_comp #(.LEN(1))
    and_comp_677 (.and_comp_in_1(w_675), .and_comp_in_2(w_676), .and_comp_out(w_677));
  or_comp #(.LEN(1))
    or_comp_678 (.or_comp_in_1(w_673), .or_comp_in_2(w_677), .or_comp_out(w_678));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_679 (.slice_in_1(w_1), .slice_out(w_679));
  eq #(.LEN(3))
    eq_680 (.eq_in_1(w_679), .eq_in_2(3'd6), .eq_out(w_680));
  and_comp #(.LEN(1))
    and_comp_681 (.and_comp_in_1(w_680), .and_comp_in_2(w_662), .and_comp_out(w_681));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_682 (.slice_in_1(w_1), .slice_out(w_682));
  eq #(.LEN(3))
    eq_683 (.eq_in_1(w_682), .eq_in_2(3'd7), .eq_out(w_683));
  not_comp #(.LEN(1))
    not_comp_684 (.not_comp_in_1(w_662), .not_comp_out(w_684));
  and_comp #(.LEN(1))
    and_comp_685 (.and_comp_in_1(w_683), .and_comp_in_2(w_684), .and_comp_out(w_685));
  or_comp #(.LEN(1))
    or_comp_686 (.or_comp_in_1(w_681), .or_comp_in_2(w_685), .or_comp_out(w_686));
  or_comp #(.LEN(1))
    or_comp_687 (.or_comp_in_1(w_678), .or_comp_in_2(w_686), .or_comp_out(w_687));
  or_comp #(.LEN(1))
    or_comp_688 (.or_comp_in_1(w_670), .or_comp_in_2(w_687), .or_comp_out(w_688));
  add #(.LEN(32))
    add_689 (.add_in_1(w_2), .add_in_2(w_595), .add_out(w_689));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_691 (.slice_in_1(w_690), .slice_out(w_691));
  add #(.LEN(32))
    add_692 (.add_in_1(w_2), .add_in_2(32'd4), .add_out(w_692));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_694 (.slice_in_1(w_693), .slice_out(w_694));
  mux21_comp #(.LEN(32))
    mux21_comp_695 (.mux21_comp_sel(w_688), .mux21_comp_in_1(w_691), .mux21_comp_in_2(w_694), .mux21_comp_out(w_695));
  add #(.LEN(32))
    add_696 (.add_in_1(w_2), .add_in_2(32'd4), .add_out(w_696));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_698 (.slice_in_1(w_697), .slice_out(w_698));
  mux21_comp #(.LEN(32))
    mux21_comp_699 (.mux21_comp_sel(w_656), .mux21_comp_in_1(w_695), .mux21_comp_in_2(w_698), .mux21_comp_out(w_699));
  mux21_comp #(.LEN(32))
    mux21_comp_700 (.mux21_comp_sel(w_649), .mux21_comp_in_1(w_654), .mux21_comp_in_2(w_699), .mux21_comp_out(w_700));
  mux21_comp #(.LEN(32))
    mux21_comp_701 (.mux21_comp_sel(w_644), .mux21_comp_in_1(w_647), .mux21_comp_in_2(w_700), .mux21_comp_out(w_701));
  mux21_comp #(.LEN(32))
    mux21_comp_702 (.mux21_comp_sel(w_639), .mux21_comp_in_1(w_642), .mux21_comp_in_2(w_701), .mux21_comp_out(w_702));
  mux21_comp #(.LEN(32))
    mux21_comp_703 (.mux21_comp_sel(w_473), .mux21_comp_in_1(w_477), .mux21_comp_in_2(w_702), .mux21_comp_out(w_703));
  mux21_comp #(.LEN(32))
    mux21_comp_704 (.mux21_comp_sel(w_634), .mux21_comp_in_1(32'd0), .mux21_comp_in_2(w_703), .mux21_comp_out(w_704));
  not_comp #(.LEN(1))
    not_comp_705 (.not_comp_in_1(w_0), .not_comp_out(w_705));
  mux21_comp #(.LEN(5))
    mux21_comp_706 (.mux21_comp_sel(w_474), .mux21_comp_in_1(5'd0), .mux21_comp_in_2(w_475), .mux21_comp_out(w_706));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_707 (.slice_in_1(w_1), .slice_out(w_707));
  eq #(.LEN(7))
    eq_708 (.eq_in_1(w_707), .eq_in_2(7'd111), .eq_out(w_708));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_709 (.slice_in_1(w_1), .slice_out(w_709));
  eq #(.LEN(7))
    eq_710 (.eq_in_1(w_709), .eq_in_2(7'd103), .eq_out(w_710));
  or_comp #(.LEN(1))
    or_comp_711 (.or_comp_in_1(w_708), .or_comp_in_2(w_710), .or_comp_out(w_711));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_712 (.slice_in_1(w_1), .slice_out(w_712));
  eq #(.LEN(7))
    eq_713 (.eq_in_1(w_712), .eq_in_2(7'd23), .eq_out(w_713));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_714 (.slice_in_1(w_1), .slice_out(w_714));
  eq #(.LEN(7))
    eq_715 (.eq_in_1(w_714), .eq_in_2(7'd55), .eq_out(w_715));
  or_comp #(.LEN(1))
    or_comp_716 (.or_comp_in_1(w_713), .or_comp_in_2(w_715), .or_comp_out(w_716));
  or_comp #(.LEN(1))
    or_comp_717 (.or_comp_in_1(w_711), .or_comp_in_2(w_716), .or_comp_out(w_717));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_718 (.slice_in_1(w_1), .slice_out(w_718));
  eq #(.LEN(7))
    eq_719 (.eq_in_1(w_718), .eq_in_2(7'd19), .eq_out(w_719));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_720 (.slice_in_1(w_1), .slice_out(w_720));
  eq #(.LEN(7))
    eq_721 (.eq_in_1(w_720), .eq_in_2(7'd51), .eq_out(w_721));
  or_comp #(.LEN(1))
    or_comp_722 (.or_comp_in_1(w_719), .or_comp_in_2(w_721), .or_comp_out(w_722));
  or_comp #(.LEN(1))
    or_comp_723 (.or_comp_in_1(w_717), .or_comp_in_2(w_722), .or_comp_out(w_723));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_724 (.slice_in_1(w_1), .slice_out(w_724));
  mux21_comp #(.LEN(5))
    mux21_comp_725 (.mux21_comp_sel(w_723), .mux21_comp_in_1(w_724), .mux21_comp_in_2(5'd0), .mux21_comp_out(w_725));
  mux21_comp #(.LEN(5))
    mux21_comp_726 (.mux21_comp_sel(w_473), .mux21_comp_in_1(w_706), .mux21_comp_in_2(w_725), .mux21_comp_out(w_726));
  mux21_comp #(.LEN(5))
    mux21_comp_727 (.mux21_comp_sel(w_705), .mux21_comp_in_1(5'd0), .mux21_comp_in_2(w_726), .mux21_comp_out(w_727));
  eq #(.LEN(3))
    eq_728 (.eq_in_1(w_478), .eq_in_2(3'd1), .eq_out(w_728));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_729 (.slice_in_1(w_1), .slice_out(w_729));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_730 (.slice_in_1(w_1), .slice_out(w_730));
  concat #(.LEN1(7), .LEN2(5))
    concat_731 (.concat_in_1(w_729), .concat_in_2(w_730), .concat_out(w_731));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_732 (.slice_in_1(w_1), .slice_out(w_732));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_733 (.slice_in_1(w_1), .slice_out(w_733));
  concat #(.LEN1(5), .LEN2(3))
    concat_734 (.concat_in_1(w_732), .concat_in_2(w_733), .concat_out(w_734));
  concat #(.LEN1(12), .LEN2(8))
    concat_735 (.concat_in_1(w_731), .concat_in_2(w_734), .concat_out(w_735));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_736 (.slice_in_1(w_1), .slice_out(w_736));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_737 (.slice_in_1(w_1), .slice_out(w_737));
  concat #(.LEN1(5), .LEN2(7))
    concat_738 (.concat_in_1(w_736), .concat_in_2(w_737), .concat_out(w_738));
  concat #(.LEN1(20), .LEN2(12))
    concat_739 (.concat_in_1(w_735), .concat_in_2(w_738), .concat_out(w_739));
  slice #(.LEN(32), .LOWER(0), .UPPER(16))
    slice_740 (.slice_in_1(w_739), .slice_out(w_740));
  slice #(.LEN(16), .LOWER(15), .UPPER(16))
    slice_741 (.slice_in_1(w_740), .slice_out(w_741));
  not_comp #(.LEN(16))
    not_comp_742 (.not_comp_in_1(16'd0), .not_comp_out(w_742));
  mux21_comp #(.LEN(16))
    mux21_comp_743 (.mux21_comp_sel(w_741), .mux21_comp_in_1(w_742), .mux21_comp_in_2(16'd0), .mux21_comp_out(w_743));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_744 (.slice_in_1(w_1), .slice_out(w_744));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_745 (.slice_in_1(w_1), .slice_out(w_745));
  concat #(.LEN1(7), .LEN2(5))
    concat_746 (.concat_in_1(w_744), .concat_in_2(w_745), .concat_out(w_746));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_747 (.slice_in_1(w_1), .slice_out(w_747));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_748 (.slice_in_1(w_1), .slice_out(w_748));
  concat #(.LEN1(5), .LEN2(3))
    concat_749 (.concat_in_1(w_747), .concat_in_2(w_748), .concat_out(w_749));
  concat #(.LEN1(12), .LEN2(8))
    concat_750 (.concat_in_1(w_746), .concat_in_2(w_749), .concat_out(w_750));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_751 (.slice_in_1(w_1), .slice_out(w_751));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_752 (.slice_in_1(w_1), .slice_out(w_752));
  concat #(.LEN1(5), .LEN2(7))
    concat_753 (.concat_in_1(w_751), .concat_in_2(w_752), .concat_out(w_753));
  concat #(.LEN1(20), .LEN2(12))
    concat_754 (.concat_in_1(w_750), .concat_in_2(w_753), .concat_out(w_754));
  slice #(.LEN(32), .LOWER(0), .UPPER(16))
    slice_755 (.slice_in_1(w_754), .slice_out(w_755));
  concat #(.LEN1(16), .LEN2(16))
    concat_756 (.concat_in_1(w_743), .concat_in_2(w_755), .concat_out(w_756));
  eq #(.LEN(3))
    eq_757 (.eq_in_1(w_478), .eq_in_2(3'd0), .eq_out(w_757));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_758 (.slice_in_1(w_1), .slice_out(w_758));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_759 (.slice_in_1(w_1), .slice_out(w_759));
  concat #(.LEN1(7), .LEN2(5))
    concat_760 (.concat_in_1(w_758), .concat_in_2(w_759), .concat_out(w_760));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_761 (.slice_in_1(w_1), .slice_out(w_761));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_762 (.slice_in_1(w_1), .slice_out(w_762));
  concat #(.LEN1(5), .LEN2(3))
    concat_763 (.concat_in_1(w_761), .concat_in_2(w_762), .concat_out(w_763));
  concat #(.LEN1(12), .LEN2(8))
    concat_764 (.concat_in_1(w_760), .concat_in_2(w_763), .concat_out(w_764));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_765 (.slice_in_1(w_1), .slice_out(w_765));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_766 (.slice_in_1(w_1), .slice_out(w_766));
  concat #(.LEN1(5), .LEN2(7))
    concat_767 (.concat_in_1(w_765), .concat_in_2(w_766), .concat_out(w_767));
  concat #(.LEN1(20), .LEN2(12))
    concat_768 (.concat_in_1(w_764), .concat_in_2(w_767), .concat_out(w_768));
  slice #(.LEN(32), .LOWER(0), .UPPER(8))
    slice_769 (.slice_in_1(w_768), .slice_out(w_769));
  slice #(.LEN(8), .LOWER(7), .UPPER(8))
    slice_770 (.slice_in_1(w_769), .slice_out(w_770));
  not_comp #(.LEN(24))
    not_comp_771 (.not_comp_in_1(24'd0), .not_comp_out(w_771));
  mux21_comp #(.LEN(24))
    mux21_comp_772 (.mux21_comp_sel(w_770), .mux21_comp_in_1(w_771), .mux21_comp_in_2(24'd0), .mux21_comp_out(w_772));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_773 (.slice_in_1(w_1), .slice_out(w_773));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_774 (.slice_in_1(w_1), .slice_out(w_774));
  concat #(.LEN1(7), .LEN2(5))
    concat_775 (.concat_in_1(w_773), .concat_in_2(w_774), .concat_out(w_775));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_776 (.slice_in_1(w_1), .slice_out(w_776));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_777 (.slice_in_1(w_1), .slice_out(w_777));
  concat #(.LEN1(5), .LEN2(3))
    concat_778 (.concat_in_1(w_776), .concat_in_2(w_777), .concat_out(w_778));
  concat #(.LEN1(12), .LEN2(8))
    concat_779 (.concat_in_1(w_775), .concat_in_2(w_778), .concat_out(w_779));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_780 (.slice_in_1(w_1), .slice_out(w_780));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_781 (.slice_in_1(w_1), .slice_out(w_781));
  concat #(.LEN1(5), .LEN2(7))
    concat_782 (.concat_in_1(w_780), .concat_in_2(w_781), .concat_out(w_782));
  concat #(.LEN1(20), .LEN2(12))
    concat_783 (.concat_in_1(w_779), .concat_in_2(w_782), .concat_out(w_783));
  slice #(.LEN(32), .LOWER(0), .UPPER(8))
    slice_784 (.slice_in_1(w_783), .slice_out(w_784));
  concat #(.LEN1(24), .LEN2(8))
    concat_785 (.concat_in_1(w_772), .concat_in_2(w_784), .concat_out(w_785));
  eq #(.LEN(3))
    eq_786 (.eq_in_1(w_478), .eq_in_2(3'd5), .eq_out(w_786));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_787 (.slice_in_1(w_1), .slice_out(w_787));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_788 (.slice_in_1(w_1), .slice_out(w_788));
  concat #(.LEN1(7), .LEN2(5))
    concat_789 (.concat_in_1(w_787), .concat_in_2(w_788), .concat_out(w_789));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_790 (.slice_in_1(w_1), .slice_out(w_790));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_791 (.slice_in_1(w_1), .slice_out(w_791));
  concat #(.LEN1(5), .LEN2(3))
    concat_792 (.concat_in_1(w_790), .concat_in_2(w_791), .concat_out(w_792));
  concat #(.LEN1(12), .LEN2(8))
    concat_793 (.concat_in_1(w_789), .concat_in_2(w_792), .concat_out(w_793));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_794 (.slice_in_1(w_1), .slice_out(w_794));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_795 (.slice_in_1(w_1), .slice_out(w_795));
  concat #(.LEN1(5), .LEN2(7))
    concat_796 (.concat_in_1(w_794), .concat_in_2(w_795), .concat_out(w_796));
  concat #(.LEN1(20), .LEN2(12))
    concat_797 (.concat_in_1(w_793), .concat_in_2(w_796), .concat_out(w_797));
  slice #(.LEN(32), .LOWER(0), .UPPER(16))
    slice_798 (.slice_in_1(w_797), .slice_out(w_798));
  concat #(.LEN1(16), .LEN2(16))
    concat_799 (.concat_in_1(16'd0), .concat_in_2(w_798), .concat_out(w_799));
  eq #(.LEN(3))
    eq_800 (.eq_in_1(w_478), .eq_in_2(3'd4), .eq_out(w_800));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_801 (.slice_in_1(w_1), .slice_out(w_801));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_802 (.slice_in_1(w_1), .slice_out(w_802));
  concat #(.LEN1(7), .LEN2(5))
    concat_803 (.concat_in_1(w_801), .concat_in_2(w_802), .concat_out(w_803));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_804 (.slice_in_1(w_1), .slice_out(w_804));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_805 (.slice_in_1(w_1), .slice_out(w_805));
  concat #(.LEN1(5), .LEN2(3))
    concat_806 (.concat_in_1(w_804), .concat_in_2(w_805), .concat_out(w_806));
  concat #(.LEN1(12), .LEN2(8))
    concat_807 (.concat_in_1(w_803), .concat_in_2(w_806), .concat_out(w_807));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_808 (.slice_in_1(w_1), .slice_out(w_808));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_809 (.slice_in_1(w_1), .slice_out(w_809));
  concat #(.LEN1(5), .LEN2(7))
    concat_810 (.concat_in_1(w_808), .concat_in_2(w_809), .concat_out(w_810));
  concat #(.LEN1(20), .LEN2(12))
    concat_811 (.concat_in_1(w_807), .concat_in_2(w_810), .concat_out(w_811));
  slice #(.LEN(32), .LOWER(0), .UPPER(8))
    slice_812 (.slice_in_1(w_811), .slice_out(w_812));
  concat #(.LEN1(24), .LEN2(8))
    concat_813 (.concat_in_1(24'd0), .concat_in_2(w_812), .concat_out(w_813));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_814 (.slice_in_1(w_1), .slice_out(w_814));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_815 (.slice_in_1(w_1), .slice_out(w_815));
  concat #(.LEN1(7), .LEN2(5))
    concat_816 (.concat_in_1(w_814), .concat_in_2(w_815), .concat_out(w_816));
  slice #(.LEN(32), .LOWER(15), .UPPER(20))
    slice_817 (.slice_in_1(w_1), .slice_out(w_817));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_818 (.slice_in_1(w_1), .slice_out(w_818));
  concat #(.LEN1(5), .LEN2(3))
    concat_819 (.concat_in_1(w_817), .concat_in_2(w_818), .concat_out(w_819));
  concat #(.LEN1(12), .LEN2(8))
    concat_820 (.concat_in_1(w_816), .concat_in_2(w_819), .concat_out(w_820));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_821 (.slice_in_1(w_1), .slice_out(w_821));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_822 (.slice_in_1(w_1), .slice_out(w_822));
  concat #(.LEN1(5), .LEN2(7))
    concat_823 (.concat_in_1(w_821), .concat_in_2(w_822), .concat_out(w_823));
  concat #(.LEN1(20), .LEN2(12))
    concat_824 (.concat_in_1(w_820), .concat_in_2(w_823), .concat_out(w_824));
  mux21_comp #(.LEN(32))
    mux21_comp_825 (.mux21_comp_sel(w_800), .mux21_comp_in_1(w_813), .mux21_comp_in_2(w_824), .mux21_comp_out(w_825));
  mux21_comp #(.LEN(32))
    mux21_comp_826 (.mux21_comp_sel(w_786), .mux21_comp_in_1(w_799), .mux21_comp_in_2(w_825), .mux21_comp_out(w_826));
  mux21_comp #(.LEN(32))
    mux21_comp_827 (.mux21_comp_sel(w_757), .mux21_comp_in_1(w_785), .mux21_comp_in_2(w_826), .mux21_comp_out(w_827));
  mux21_comp #(.LEN(32))
    mux21_comp_828 (.mux21_comp_sel(w_728), .mux21_comp_in_1(w_756), .mux21_comp_in_2(w_827), .mux21_comp_out(w_828));
  mux21_comp #(.LEN(32))
    mux21_comp_829 (.mux21_comp_sel(w_474), .mux21_comp_in_1(32'd0), .mux21_comp_in_2(w_828), .mux21_comp_out(w_829));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_830 (.slice_in_1(w_1), .slice_out(w_830));
  eq #(.LEN(7))
    eq_831 (.eq_in_1(w_830), .eq_in_2(7'd55), .eq_out(w_831));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_832 (.slice_in_1(w_1), .slice_out(w_832));
  eq #(.LEN(7))
    eq_833 (.eq_in_1(w_832), .eq_in_2(7'd23), .eq_out(w_833));
  add #(.LEN(32))
    add_834 (.add_in_1(w_2), .add_in_2(w_595), .add_out(w_834));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_836 (.slice_in_1(w_835), .slice_out(w_836));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_837 (.slice_in_1(w_1), .slice_out(w_837));
  eq #(.LEN(7))
    eq_838 (.eq_in_1(w_837), .eq_in_2(7'd111), .eq_out(w_838));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_839 (.slice_in_1(w_1), .slice_out(w_839));
  eq #(.LEN(7))
    eq_840 (.eq_in_1(w_839), .eq_in_2(7'd103), .eq_out(w_840));
  or_comp #(.LEN(1))
    or_comp_841 (.or_comp_in_1(w_838), .or_comp_in_2(w_840), .or_comp_out(w_841));
  add #(.LEN(32))
    add_842 (.add_in_1(w_2), .add_in_2(32'd4), .add_out(w_842));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_844 (.slice_in_1(w_843), .slice_out(w_844));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_845 (.slice_in_1(w_1), .slice_out(w_845));
  eq #(.LEN(7))
    eq_846 (.eq_in_1(w_845), .eq_in_2(7'd51), .eq_out(w_846));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_847 (.slice_in_1(w_1), .slice_out(w_847));
  eq #(.LEN(7))
    eq_848 (.eq_in_1(w_847), .eq_in_2(7'd19), .eq_out(w_848));
  or_comp #(.LEN(1))
    or_comp_849 (.or_comp_in_1(w_846), .or_comp_in_2(w_848), .or_comp_out(w_849));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_850 (.slice_in_1(w_1), .slice_out(w_850));
  eq #(.LEN(3))
    eq_851 (.eq_in_1(w_850), .eq_in_2(3'd0), .eq_out(w_851));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_852 (.slice_in_1(w_1), .slice_out(w_852));
  eq #(.LEN(7))
    eq_853 (.eq_in_1(w_852), .eq_in_2(7'd19), .eq_out(w_853));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_854 (.slice_in_1(w_1), .slice_out(w_854));
  eq #(.LEN(7))
    eq_855 (.eq_in_1(w_854), .eq_in_2(7'd32), .eq_out(w_855));
  mux21_comp #(.LEN(10))
    mux21_comp_856 (.mux21_comp_sel(w_855), .mux21_comp_in_1(10'd2), .mux21_comp_in_2(10'd1), .mux21_comp_out(w_856));
  mux21_comp #(.LEN(10))
    mux21_comp_857 (.mux21_comp_sel(w_853), .mux21_comp_in_1(10'd1), .mux21_comp_in_2(w_856), .mux21_comp_out(w_857));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_858 (.slice_in_1(w_1), .slice_out(w_858));
  eq #(.LEN(3))
    eq_859 (.eq_in_1(w_858), .eq_in_2(3'd1), .eq_out(w_859));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_860 (.slice_in_1(w_1), .slice_out(w_860));
  eq #(.LEN(3))
    eq_861 (.eq_in_1(w_860), .eq_in_2(3'd2), .eq_out(w_861));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_862 (.slice_in_1(w_1), .slice_out(w_862));
  eq #(.LEN(3))
    eq_863 (.eq_in_1(w_862), .eq_in_2(3'd3), .eq_out(w_863));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_864 (.slice_in_1(w_1), .slice_out(w_864));
  eq #(.LEN(3))
    eq_865 (.eq_in_1(w_864), .eq_in_2(3'd4), .eq_out(w_865));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_866 (.slice_in_1(w_1), .slice_out(w_866));
  eq #(.LEN(3))
    eq_867 (.eq_in_1(w_866), .eq_in_2(3'd5), .eq_out(w_867));
  slice #(.LEN(32), .LOWER(25), .UPPER(32))
    slice_868 (.slice_in_1(w_1), .slice_out(w_868));
  eq #(.LEN(7))
    eq_869 (.eq_in_1(w_868), .eq_in_2(7'd32), .eq_out(w_869));
  mux21_comp #(.LEN(10))
    mux21_comp_870 (.mux21_comp_sel(w_869), .mux21_comp_in_1(10'd128), .mux21_comp_in_2(10'd64), .mux21_comp_out(w_870));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_871 (.slice_in_1(w_1), .slice_out(w_871));
  eq #(.LEN(3))
    eq_872 (.eq_in_1(w_871), .eq_in_2(3'd6), .eq_out(w_872));
  mux21_comp #(.LEN(10))
    mux21_comp_873 (.mux21_comp_sel(w_872), .mux21_comp_in_1(10'd256), .mux21_comp_in_2(10'd512), .mux21_comp_out(w_873));
  mux21_comp #(.LEN(10))
    mux21_comp_874 (.mux21_comp_sel(w_867), .mux21_comp_in_1(w_870), .mux21_comp_in_2(w_873), .mux21_comp_out(w_874));
  mux21_comp #(.LEN(10))
    mux21_comp_875 (.mux21_comp_sel(w_865), .mux21_comp_in_1(10'd16), .mux21_comp_in_2(w_874), .mux21_comp_out(w_875));
  mux21_comp #(.LEN(10))
    mux21_comp_876 (.mux21_comp_sel(w_863), .mux21_comp_in_1(10'd8), .mux21_comp_in_2(w_875), .mux21_comp_out(w_876));
  mux21_comp #(.LEN(10))
    mux21_comp_877 (.mux21_comp_sel(w_861), .mux21_comp_in_1(10'd4), .mux21_comp_in_2(w_876), .mux21_comp_out(w_877));
  mux21_comp #(.LEN(10))
    mux21_comp_878 (.mux21_comp_sel(w_859), .mux21_comp_in_1(10'd32), .mux21_comp_in_2(w_877), .mux21_comp_out(w_878));
  mux21_comp #(.LEN(10))
    mux21_comp_879 (.mux21_comp_sel(w_851), .mux21_comp_in_1(w_857), .mux21_comp_in_2(w_878), .mux21_comp_out(w_879));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_880 (.slice_in_1(w_1), .slice_out(w_880));
  eq #(.LEN(7))
    eq_881 (.eq_in_1(w_880), .eq_in_2(7'd51), .eq_out(w_881));
  mux21_comp #(.LEN(32))
    mux21_comp_882 (.mux21_comp_sel(w_881), .mux21_comp_in_1(w_472), .mux21_comp_in_2(w_595), .mux21_comp_out(w_882));
  slice #(.LEN(10), .LOWER(0), .UPPER(1))
    slice_886 (.slice_in_1(w_883), .slice_out(w_886));
  add #(.LEN(32))
    add_887 (.add_in_1(w_884), .add_in_2(w_885), .add_out(w_887));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_889 (.slice_in_1(w_888), .slice_out(w_889));
  slice #(.LEN(10), .LOWER(1), .UPPER(2))
    slice_890 (.slice_in_1(w_883), .slice_out(w_890));
  not_comp #(.LEN(32))
    not_comp_891 (.not_comp_in_1(w_885), .not_comp_out(w_891));
  add #(.LEN(32))
    add_892 (.add_in_1(w_891), .add_in_2(32'd1), .add_out(w_892));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_894 (.slice_in_1(w_893), .slice_out(w_894));
  add #(.LEN(32))
    add_895 (.add_in_1(w_884), .add_in_2(w_894), .add_out(w_895));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_897 (.slice_in_1(w_896), .slice_out(w_897));
  slice #(.LEN(10), .LOWER(2), .UPPER(3))
    slice_898 (.slice_in_1(w_883), .slice_out(w_898));
  lt #(.LEN(32))
    lt_899 (.lt_in_1(w_884), .lt_in_2(w_885), .lt_out(w_899));
  mux21_comp #(.LEN(32))
    mux21_comp_900 (.mux21_comp_sel(w_899), .mux21_comp_in_1(32'd1), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_900));
  slice #(.LEN(10), .LOWER(3), .UPPER(4))
    slice_901 (.slice_in_1(w_883), .slice_out(w_901));
  ltu #(.LEN(32))
    ltu_902 (.ltu_in_1(w_884), .ltu_in_2(w_885), .ltu_out(w_902));
  mux21_comp #(.LEN(32))
    mux21_comp_903 (.mux21_comp_sel(w_902), .mux21_comp_in_1(32'd1), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_903));
  slice #(.LEN(10), .LOWER(4), .UPPER(5))
    slice_904 (.slice_in_1(w_883), .slice_out(w_904));
  xor_comp #(.LEN(32))
    xor_comp_905 (.xor_comp_in_1(w_884), .xor_comp_in_2(w_885), .xor_comp_out(w_905));
  slice #(.LEN(10), .LOWER(5), .UPPER(6))
    slice_906 (.slice_in_1(w_883), .slice_out(w_906));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_907 (.slice_in_1(w_885), .slice_out(w_907));
  eq #(.LEN(5))
    eq_908 (.eq_in_1(w_907), .eq_in_2(5'd31), .eq_out(w_908));
  sll #(.LEN(32), .SHAMT(31))
    sll_909 (.sll_in_1(w_884), .sll_out(w_909));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_910 (.slice_in_1(w_885), .slice_out(w_910));
  eq #(.LEN(5))
    eq_911 (.eq_in_1(w_910), .eq_in_2(5'd30), .eq_out(w_911));
  sll #(.LEN(32), .SHAMT(30))
    sll_912 (.sll_in_1(w_884), .sll_out(w_912));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_913 (.slice_in_1(w_885), .slice_out(w_913));
  eq #(.LEN(5))
    eq_914 (.eq_in_1(w_913), .eq_in_2(5'd29), .eq_out(w_914));
  sll #(.LEN(32), .SHAMT(29))
    sll_915 (.sll_in_1(w_884), .sll_out(w_915));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_916 (.slice_in_1(w_885), .slice_out(w_916));
  eq #(.LEN(5))
    eq_917 (.eq_in_1(w_916), .eq_in_2(5'd28), .eq_out(w_917));
  sll #(.LEN(32), .SHAMT(28))
    sll_918 (.sll_in_1(w_884), .sll_out(w_918));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_919 (.slice_in_1(w_885), .slice_out(w_919));
  eq #(.LEN(5))
    eq_920 (.eq_in_1(w_919), .eq_in_2(5'd27), .eq_out(w_920));
  sll #(.LEN(32), .SHAMT(27))
    sll_921 (.sll_in_1(w_884), .sll_out(w_921));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_922 (.slice_in_1(w_885), .slice_out(w_922));
  eq #(.LEN(5))
    eq_923 (.eq_in_1(w_922), .eq_in_2(5'd26), .eq_out(w_923));
  sll #(.LEN(32), .SHAMT(26))
    sll_924 (.sll_in_1(w_884), .sll_out(w_924));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_925 (.slice_in_1(w_885), .slice_out(w_925));
  eq #(.LEN(5))
    eq_926 (.eq_in_1(w_925), .eq_in_2(5'd25), .eq_out(w_926));
  sll #(.LEN(32), .SHAMT(25))
    sll_927 (.sll_in_1(w_884), .sll_out(w_927));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_928 (.slice_in_1(w_885), .slice_out(w_928));
  eq #(.LEN(5))
    eq_929 (.eq_in_1(w_928), .eq_in_2(5'd24), .eq_out(w_929));
  sll #(.LEN(32), .SHAMT(24))
    sll_930 (.sll_in_1(w_884), .sll_out(w_930));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_931 (.slice_in_1(w_885), .slice_out(w_931));
  eq #(.LEN(5))
    eq_932 (.eq_in_1(w_931), .eq_in_2(5'd23), .eq_out(w_932));
  sll #(.LEN(32), .SHAMT(23))
    sll_933 (.sll_in_1(w_884), .sll_out(w_933));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_934 (.slice_in_1(w_885), .slice_out(w_934));
  eq #(.LEN(5))
    eq_935 (.eq_in_1(w_934), .eq_in_2(5'd22), .eq_out(w_935));
  sll #(.LEN(32), .SHAMT(22))
    sll_936 (.sll_in_1(w_884), .sll_out(w_936));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_937 (.slice_in_1(w_885), .slice_out(w_937));
  eq #(.LEN(5))
    eq_938 (.eq_in_1(w_937), .eq_in_2(5'd21), .eq_out(w_938));
  sll #(.LEN(32), .SHAMT(21))
    sll_939 (.sll_in_1(w_884), .sll_out(w_939));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_940 (.slice_in_1(w_885), .slice_out(w_940));
  eq #(.LEN(5))
    eq_941 (.eq_in_1(w_940), .eq_in_2(5'd20), .eq_out(w_941));
  sll #(.LEN(32), .SHAMT(20))
    sll_942 (.sll_in_1(w_884), .sll_out(w_942));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_943 (.slice_in_1(w_885), .slice_out(w_943));
  eq #(.LEN(5))
    eq_944 (.eq_in_1(w_943), .eq_in_2(5'd19), .eq_out(w_944));
  sll #(.LEN(32), .SHAMT(19))
    sll_945 (.sll_in_1(w_884), .sll_out(w_945));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_946 (.slice_in_1(w_885), .slice_out(w_946));
  eq #(.LEN(5))
    eq_947 (.eq_in_1(w_946), .eq_in_2(5'd18), .eq_out(w_947));
  sll #(.LEN(32), .SHAMT(18))
    sll_948 (.sll_in_1(w_884), .sll_out(w_948));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_949 (.slice_in_1(w_885), .slice_out(w_949));
  eq #(.LEN(5))
    eq_950 (.eq_in_1(w_949), .eq_in_2(5'd17), .eq_out(w_950));
  sll #(.LEN(32), .SHAMT(17))
    sll_951 (.sll_in_1(w_884), .sll_out(w_951));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_952 (.slice_in_1(w_885), .slice_out(w_952));
  eq #(.LEN(5))
    eq_953 (.eq_in_1(w_952), .eq_in_2(5'd16), .eq_out(w_953));
  sll #(.LEN(32), .SHAMT(16))
    sll_954 (.sll_in_1(w_884), .sll_out(w_954));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_955 (.slice_in_1(w_885), .slice_out(w_955));
  eq #(.LEN(5))
    eq_956 (.eq_in_1(w_955), .eq_in_2(5'd15), .eq_out(w_956));
  sll #(.LEN(32), .SHAMT(15))
    sll_957 (.sll_in_1(w_884), .sll_out(w_957));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_958 (.slice_in_1(w_885), .slice_out(w_958));
  eq #(.LEN(5))
    eq_959 (.eq_in_1(w_958), .eq_in_2(5'd14), .eq_out(w_959));
  sll #(.LEN(32), .SHAMT(14))
    sll_960 (.sll_in_1(w_884), .sll_out(w_960));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_961 (.slice_in_1(w_885), .slice_out(w_961));
  eq #(.LEN(5))
    eq_962 (.eq_in_1(w_961), .eq_in_2(5'd13), .eq_out(w_962));
  sll #(.LEN(32), .SHAMT(13))
    sll_963 (.sll_in_1(w_884), .sll_out(w_963));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_964 (.slice_in_1(w_885), .slice_out(w_964));
  eq #(.LEN(5))
    eq_965 (.eq_in_1(w_964), .eq_in_2(5'd12), .eq_out(w_965));
  sll #(.LEN(32), .SHAMT(12))
    sll_966 (.sll_in_1(w_884), .sll_out(w_966));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_967 (.slice_in_1(w_885), .slice_out(w_967));
  eq #(.LEN(5))
    eq_968 (.eq_in_1(w_967), .eq_in_2(5'd11), .eq_out(w_968));
  sll #(.LEN(32), .SHAMT(11))
    sll_969 (.sll_in_1(w_884), .sll_out(w_969));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_970 (.slice_in_1(w_885), .slice_out(w_970));
  eq #(.LEN(5))
    eq_971 (.eq_in_1(w_970), .eq_in_2(5'd10), .eq_out(w_971));
  sll #(.LEN(32), .SHAMT(10))
    sll_972 (.sll_in_1(w_884), .sll_out(w_972));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_973 (.slice_in_1(w_885), .slice_out(w_973));
  eq #(.LEN(5))
    eq_974 (.eq_in_1(w_973), .eq_in_2(5'd9), .eq_out(w_974));
  sll #(.LEN(32), .SHAMT(9))
    sll_975 (.sll_in_1(w_884), .sll_out(w_975));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_976 (.slice_in_1(w_885), .slice_out(w_976));
  eq #(.LEN(5))
    eq_977 (.eq_in_1(w_976), .eq_in_2(5'd8), .eq_out(w_977));
  sll #(.LEN(32), .SHAMT(8))
    sll_978 (.sll_in_1(w_884), .sll_out(w_978));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_979 (.slice_in_1(w_885), .slice_out(w_979));
  eq #(.LEN(5))
    eq_980 (.eq_in_1(w_979), .eq_in_2(5'd7), .eq_out(w_980));
  sll #(.LEN(32), .SHAMT(7))
    sll_981 (.sll_in_1(w_884), .sll_out(w_981));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_982 (.slice_in_1(w_885), .slice_out(w_982));
  eq #(.LEN(5))
    eq_983 (.eq_in_1(w_982), .eq_in_2(5'd6), .eq_out(w_983));
  sll #(.LEN(32), .SHAMT(6))
    sll_984 (.sll_in_1(w_884), .sll_out(w_984));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_985 (.slice_in_1(w_885), .slice_out(w_985));
  eq #(.LEN(5))
    eq_986 (.eq_in_1(w_985), .eq_in_2(5'd5), .eq_out(w_986));
  sll #(.LEN(32), .SHAMT(5))
    sll_987 (.sll_in_1(w_884), .sll_out(w_987));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_988 (.slice_in_1(w_885), .slice_out(w_988));
  eq #(.LEN(5))
    eq_989 (.eq_in_1(w_988), .eq_in_2(5'd4), .eq_out(w_989));
  sll #(.LEN(32), .SHAMT(4))
    sll_990 (.sll_in_1(w_884), .sll_out(w_990));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_991 (.slice_in_1(w_885), .slice_out(w_991));
  eq #(.LEN(5))
    eq_992 (.eq_in_1(w_991), .eq_in_2(5'd3), .eq_out(w_992));
  sll #(.LEN(32), .SHAMT(3))
    sll_993 (.sll_in_1(w_884), .sll_out(w_993));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_994 (.slice_in_1(w_885), .slice_out(w_994));
  eq #(.LEN(5))
    eq_995 (.eq_in_1(w_994), .eq_in_2(5'd2), .eq_out(w_995));
  sll #(.LEN(32), .SHAMT(2))
    sll_996 (.sll_in_1(w_884), .sll_out(w_996));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_997 (.slice_in_1(w_885), .slice_out(w_997));
  eq #(.LEN(5))
    eq_998 (.eq_in_1(w_997), .eq_in_2(5'd1), .eq_out(w_998));
  sll #(.LEN(32), .SHAMT(1))
    sll_999 (.sll_in_1(w_884), .sll_out(w_999));
  mux21_comp #(.LEN(32))
    mux21_comp_1000 (.mux21_comp_sel(w_998), .mux21_comp_in_1(w_999), .mux21_comp_in_2(w_884), .mux21_comp_out(w_1000));
  mux21_comp #(.LEN(32))
    mux21_comp_1001 (.mux21_comp_sel(w_995), .mux21_comp_in_1(w_996), .mux21_comp_in_2(w_1000), .mux21_comp_out(w_1001));
  mux21_comp #(.LEN(32))
    mux21_comp_1002 (.mux21_comp_sel(w_992), .mux21_comp_in_1(w_993), .mux21_comp_in_2(w_1001), .mux21_comp_out(w_1002));
  mux21_comp #(.LEN(32))
    mux21_comp_1003 (.mux21_comp_sel(w_989), .mux21_comp_in_1(w_990), .mux21_comp_in_2(w_1002), .mux21_comp_out(w_1003));
  mux21_comp #(.LEN(32))
    mux21_comp_1004 (.mux21_comp_sel(w_986), .mux21_comp_in_1(w_987), .mux21_comp_in_2(w_1003), .mux21_comp_out(w_1004));
  mux21_comp #(.LEN(32))
    mux21_comp_1005 (.mux21_comp_sel(w_983), .mux21_comp_in_1(w_984), .mux21_comp_in_2(w_1004), .mux21_comp_out(w_1005));
  mux21_comp #(.LEN(32))
    mux21_comp_1006 (.mux21_comp_sel(w_980), .mux21_comp_in_1(w_981), .mux21_comp_in_2(w_1005), .mux21_comp_out(w_1006));
  mux21_comp #(.LEN(32))
    mux21_comp_1007 (.mux21_comp_sel(w_977), .mux21_comp_in_1(w_978), .mux21_comp_in_2(w_1006), .mux21_comp_out(w_1007));
  mux21_comp #(.LEN(32))
    mux21_comp_1008 (.mux21_comp_sel(w_974), .mux21_comp_in_1(w_975), .mux21_comp_in_2(w_1007), .mux21_comp_out(w_1008));
  mux21_comp #(.LEN(32))
    mux21_comp_1009 (.mux21_comp_sel(w_971), .mux21_comp_in_1(w_972), .mux21_comp_in_2(w_1008), .mux21_comp_out(w_1009));
  mux21_comp #(.LEN(32))
    mux21_comp_1010 (.mux21_comp_sel(w_968), .mux21_comp_in_1(w_969), .mux21_comp_in_2(w_1009), .mux21_comp_out(w_1010));
  mux21_comp #(.LEN(32))
    mux21_comp_1011 (.mux21_comp_sel(w_965), .mux21_comp_in_1(w_966), .mux21_comp_in_2(w_1010), .mux21_comp_out(w_1011));
  mux21_comp #(.LEN(32))
    mux21_comp_1012 (.mux21_comp_sel(w_962), .mux21_comp_in_1(w_963), .mux21_comp_in_2(w_1011), .mux21_comp_out(w_1012));
  mux21_comp #(.LEN(32))
    mux21_comp_1013 (.mux21_comp_sel(w_959), .mux21_comp_in_1(w_960), .mux21_comp_in_2(w_1012), .mux21_comp_out(w_1013));
  mux21_comp #(.LEN(32))
    mux21_comp_1014 (.mux21_comp_sel(w_956), .mux21_comp_in_1(w_957), .mux21_comp_in_2(w_1013), .mux21_comp_out(w_1014));
  mux21_comp #(.LEN(32))
    mux21_comp_1015 (.mux21_comp_sel(w_953), .mux21_comp_in_1(w_954), .mux21_comp_in_2(w_1014), .mux21_comp_out(w_1015));
  mux21_comp #(.LEN(32))
    mux21_comp_1016 (.mux21_comp_sel(w_950), .mux21_comp_in_1(w_951), .mux21_comp_in_2(w_1015), .mux21_comp_out(w_1016));
  mux21_comp #(.LEN(32))
    mux21_comp_1017 (.mux21_comp_sel(w_947), .mux21_comp_in_1(w_948), .mux21_comp_in_2(w_1016), .mux21_comp_out(w_1017));
  mux21_comp #(.LEN(32))
    mux21_comp_1018 (.mux21_comp_sel(w_944), .mux21_comp_in_1(w_945), .mux21_comp_in_2(w_1017), .mux21_comp_out(w_1018));
  mux21_comp #(.LEN(32))
    mux21_comp_1019 (.mux21_comp_sel(w_941), .mux21_comp_in_1(w_942), .mux21_comp_in_2(w_1018), .mux21_comp_out(w_1019));
  mux21_comp #(.LEN(32))
    mux21_comp_1020 (.mux21_comp_sel(w_938), .mux21_comp_in_1(w_939), .mux21_comp_in_2(w_1019), .mux21_comp_out(w_1020));
  mux21_comp #(.LEN(32))
    mux21_comp_1021 (.mux21_comp_sel(w_935), .mux21_comp_in_1(w_936), .mux21_comp_in_2(w_1020), .mux21_comp_out(w_1021));
  mux21_comp #(.LEN(32))
    mux21_comp_1022 (.mux21_comp_sel(w_932), .mux21_comp_in_1(w_933), .mux21_comp_in_2(w_1021), .mux21_comp_out(w_1022));
  mux21_comp #(.LEN(32))
    mux21_comp_1023 (.mux21_comp_sel(w_929), .mux21_comp_in_1(w_930), .mux21_comp_in_2(w_1022), .mux21_comp_out(w_1023));
  mux21_comp #(.LEN(32))
    mux21_comp_1024 (.mux21_comp_sel(w_926), .mux21_comp_in_1(w_927), .mux21_comp_in_2(w_1023), .mux21_comp_out(w_1024));
  mux21_comp #(.LEN(32))
    mux21_comp_1025 (.mux21_comp_sel(w_923), .mux21_comp_in_1(w_924), .mux21_comp_in_2(w_1024), .mux21_comp_out(w_1025));
  mux21_comp #(.LEN(32))
    mux21_comp_1026 (.mux21_comp_sel(w_920), .mux21_comp_in_1(w_921), .mux21_comp_in_2(w_1025), .mux21_comp_out(w_1026));
  mux21_comp #(.LEN(32))
    mux21_comp_1027 (.mux21_comp_sel(w_917), .mux21_comp_in_1(w_918), .mux21_comp_in_2(w_1026), .mux21_comp_out(w_1027));
  mux21_comp #(.LEN(32))
    mux21_comp_1028 (.mux21_comp_sel(w_914), .mux21_comp_in_1(w_915), .mux21_comp_in_2(w_1027), .mux21_comp_out(w_1028));
  mux21_comp #(.LEN(32))
    mux21_comp_1029 (.mux21_comp_sel(w_911), .mux21_comp_in_1(w_912), .mux21_comp_in_2(w_1028), .mux21_comp_out(w_1029));
  mux21_comp #(.LEN(32))
    mux21_comp_1030 (.mux21_comp_sel(w_908), .mux21_comp_in_1(w_909), .mux21_comp_in_2(w_1029), .mux21_comp_out(w_1030));
  slice #(.LEN(10), .LOWER(6), .UPPER(7))
    slice_1031 (.slice_in_1(w_883), .slice_out(w_1031));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1032 (.slice_in_1(w_885), .slice_out(w_1032));
  eq #(.LEN(5))
    eq_1033 (.eq_in_1(w_1032), .eq_in_2(5'd31), .eq_out(w_1033));
  srl #(.LEN(32), .SHAMT(31))
    srl_1034 (.srl_in_1(w_884), .srl_out(w_1034));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1035 (.slice_in_1(w_885), .slice_out(w_1035));
  eq #(.LEN(5))
    eq_1036 (.eq_in_1(w_1035), .eq_in_2(5'd30), .eq_out(w_1036));
  srl #(.LEN(32), .SHAMT(30))
    srl_1037 (.srl_in_1(w_884), .srl_out(w_1037));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1038 (.slice_in_1(w_885), .slice_out(w_1038));
  eq #(.LEN(5))
    eq_1039 (.eq_in_1(w_1038), .eq_in_2(5'd29), .eq_out(w_1039));
  srl #(.LEN(32), .SHAMT(29))
    srl_1040 (.srl_in_1(w_884), .srl_out(w_1040));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1041 (.slice_in_1(w_885), .slice_out(w_1041));
  eq #(.LEN(5))
    eq_1042 (.eq_in_1(w_1041), .eq_in_2(5'd28), .eq_out(w_1042));
  srl #(.LEN(32), .SHAMT(28))
    srl_1043 (.srl_in_1(w_884), .srl_out(w_1043));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1044 (.slice_in_1(w_885), .slice_out(w_1044));
  eq #(.LEN(5))
    eq_1045 (.eq_in_1(w_1044), .eq_in_2(5'd27), .eq_out(w_1045));
  srl #(.LEN(32), .SHAMT(27))
    srl_1046 (.srl_in_1(w_884), .srl_out(w_1046));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1047 (.slice_in_1(w_885), .slice_out(w_1047));
  eq #(.LEN(5))
    eq_1048 (.eq_in_1(w_1047), .eq_in_2(5'd26), .eq_out(w_1048));
  srl #(.LEN(32), .SHAMT(26))
    srl_1049 (.srl_in_1(w_884), .srl_out(w_1049));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1050 (.slice_in_1(w_885), .slice_out(w_1050));
  eq #(.LEN(5))
    eq_1051 (.eq_in_1(w_1050), .eq_in_2(5'd25), .eq_out(w_1051));
  srl #(.LEN(32), .SHAMT(25))
    srl_1052 (.srl_in_1(w_884), .srl_out(w_1052));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1053 (.slice_in_1(w_885), .slice_out(w_1053));
  eq #(.LEN(5))
    eq_1054 (.eq_in_1(w_1053), .eq_in_2(5'd24), .eq_out(w_1054));
  srl #(.LEN(32), .SHAMT(24))
    srl_1055 (.srl_in_1(w_884), .srl_out(w_1055));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1056 (.slice_in_1(w_885), .slice_out(w_1056));
  eq #(.LEN(5))
    eq_1057 (.eq_in_1(w_1056), .eq_in_2(5'd23), .eq_out(w_1057));
  srl #(.LEN(32), .SHAMT(23))
    srl_1058 (.srl_in_1(w_884), .srl_out(w_1058));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1059 (.slice_in_1(w_885), .slice_out(w_1059));
  eq #(.LEN(5))
    eq_1060 (.eq_in_1(w_1059), .eq_in_2(5'd22), .eq_out(w_1060));
  srl #(.LEN(32), .SHAMT(22))
    srl_1061 (.srl_in_1(w_884), .srl_out(w_1061));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1062 (.slice_in_1(w_885), .slice_out(w_1062));
  eq #(.LEN(5))
    eq_1063 (.eq_in_1(w_1062), .eq_in_2(5'd21), .eq_out(w_1063));
  srl #(.LEN(32), .SHAMT(21))
    srl_1064 (.srl_in_1(w_884), .srl_out(w_1064));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1065 (.slice_in_1(w_885), .slice_out(w_1065));
  eq #(.LEN(5))
    eq_1066 (.eq_in_1(w_1065), .eq_in_2(5'd20), .eq_out(w_1066));
  srl #(.LEN(32), .SHAMT(20))
    srl_1067 (.srl_in_1(w_884), .srl_out(w_1067));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1068 (.slice_in_1(w_885), .slice_out(w_1068));
  eq #(.LEN(5))
    eq_1069 (.eq_in_1(w_1068), .eq_in_2(5'd19), .eq_out(w_1069));
  srl #(.LEN(32), .SHAMT(19))
    srl_1070 (.srl_in_1(w_884), .srl_out(w_1070));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1071 (.slice_in_1(w_885), .slice_out(w_1071));
  eq #(.LEN(5))
    eq_1072 (.eq_in_1(w_1071), .eq_in_2(5'd18), .eq_out(w_1072));
  srl #(.LEN(32), .SHAMT(18))
    srl_1073 (.srl_in_1(w_884), .srl_out(w_1073));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1074 (.slice_in_1(w_885), .slice_out(w_1074));
  eq #(.LEN(5))
    eq_1075 (.eq_in_1(w_1074), .eq_in_2(5'd17), .eq_out(w_1075));
  srl #(.LEN(32), .SHAMT(17))
    srl_1076 (.srl_in_1(w_884), .srl_out(w_1076));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1077 (.slice_in_1(w_885), .slice_out(w_1077));
  eq #(.LEN(5))
    eq_1078 (.eq_in_1(w_1077), .eq_in_2(5'd16), .eq_out(w_1078));
  srl #(.LEN(32), .SHAMT(16))
    srl_1079 (.srl_in_1(w_884), .srl_out(w_1079));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1080 (.slice_in_1(w_885), .slice_out(w_1080));
  eq #(.LEN(5))
    eq_1081 (.eq_in_1(w_1080), .eq_in_2(5'd15), .eq_out(w_1081));
  srl #(.LEN(32), .SHAMT(15))
    srl_1082 (.srl_in_1(w_884), .srl_out(w_1082));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1083 (.slice_in_1(w_885), .slice_out(w_1083));
  eq #(.LEN(5))
    eq_1084 (.eq_in_1(w_1083), .eq_in_2(5'd14), .eq_out(w_1084));
  srl #(.LEN(32), .SHAMT(14))
    srl_1085 (.srl_in_1(w_884), .srl_out(w_1085));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1086 (.slice_in_1(w_885), .slice_out(w_1086));
  eq #(.LEN(5))
    eq_1087 (.eq_in_1(w_1086), .eq_in_2(5'd13), .eq_out(w_1087));
  srl #(.LEN(32), .SHAMT(13))
    srl_1088 (.srl_in_1(w_884), .srl_out(w_1088));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1089 (.slice_in_1(w_885), .slice_out(w_1089));
  eq #(.LEN(5))
    eq_1090 (.eq_in_1(w_1089), .eq_in_2(5'd12), .eq_out(w_1090));
  srl #(.LEN(32), .SHAMT(12))
    srl_1091 (.srl_in_1(w_884), .srl_out(w_1091));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1092 (.slice_in_1(w_885), .slice_out(w_1092));
  eq #(.LEN(5))
    eq_1093 (.eq_in_1(w_1092), .eq_in_2(5'd11), .eq_out(w_1093));
  srl #(.LEN(32), .SHAMT(11))
    srl_1094 (.srl_in_1(w_884), .srl_out(w_1094));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1095 (.slice_in_1(w_885), .slice_out(w_1095));
  eq #(.LEN(5))
    eq_1096 (.eq_in_1(w_1095), .eq_in_2(5'd10), .eq_out(w_1096));
  srl #(.LEN(32), .SHAMT(10))
    srl_1097 (.srl_in_1(w_884), .srl_out(w_1097));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1098 (.slice_in_1(w_885), .slice_out(w_1098));
  eq #(.LEN(5))
    eq_1099 (.eq_in_1(w_1098), .eq_in_2(5'd9), .eq_out(w_1099));
  srl #(.LEN(32), .SHAMT(9))
    srl_1100 (.srl_in_1(w_884), .srl_out(w_1100));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1101 (.slice_in_1(w_885), .slice_out(w_1101));
  eq #(.LEN(5))
    eq_1102 (.eq_in_1(w_1101), .eq_in_2(5'd8), .eq_out(w_1102));
  srl #(.LEN(32), .SHAMT(8))
    srl_1103 (.srl_in_1(w_884), .srl_out(w_1103));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1104 (.slice_in_1(w_885), .slice_out(w_1104));
  eq #(.LEN(5))
    eq_1105 (.eq_in_1(w_1104), .eq_in_2(5'd7), .eq_out(w_1105));
  srl #(.LEN(32), .SHAMT(7))
    srl_1106 (.srl_in_1(w_884), .srl_out(w_1106));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1107 (.slice_in_1(w_885), .slice_out(w_1107));
  eq #(.LEN(5))
    eq_1108 (.eq_in_1(w_1107), .eq_in_2(5'd6), .eq_out(w_1108));
  srl #(.LEN(32), .SHAMT(6))
    srl_1109 (.srl_in_1(w_884), .srl_out(w_1109));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1110 (.slice_in_1(w_885), .slice_out(w_1110));
  eq #(.LEN(5))
    eq_1111 (.eq_in_1(w_1110), .eq_in_2(5'd5), .eq_out(w_1111));
  srl #(.LEN(32), .SHAMT(5))
    srl_1112 (.srl_in_1(w_884), .srl_out(w_1112));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1113 (.slice_in_1(w_885), .slice_out(w_1113));
  eq #(.LEN(5))
    eq_1114 (.eq_in_1(w_1113), .eq_in_2(5'd4), .eq_out(w_1114));
  srl #(.LEN(32), .SHAMT(4))
    srl_1115 (.srl_in_1(w_884), .srl_out(w_1115));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1116 (.slice_in_1(w_885), .slice_out(w_1116));
  eq #(.LEN(5))
    eq_1117 (.eq_in_1(w_1116), .eq_in_2(5'd3), .eq_out(w_1117));
  srl #(.LEN(32), .SHAMT(3))
    srl_1118 (.srl_in_1(w_884), .srl_out(w_1118));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1119 (.slice_in_1(w_885), .slice_out(w_1119));
  eq #(.LEN(5))
    eq_1120 (.eq_in_1(w_1119), .eq_in_2(5'd2), .eq_out(w_1120));
  srl #(.LEN(32), .SHAMT(2))
    srl_1121 (.srl_in_1(w_884), .srl_out(w_1121));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1122 (.slice_in_1(w_885), .slice_out(w_1122));
  eq #(.LEN(5))
    eq_1123 (.eq_in_1(w_1122), .eq_in_2(5'd1), .eq_out(w_1123));
  srl #(.LEN(32), .SHAMT(1))
    srl_1124 (.srl_in_1(w_884), .srl_out(w_1124));
  mux21_comp #(.LEN(32))
    mux21_comp_1125 (.mux21_comp_sel(w_1123), .mux21_comp_in_1(w_1124), .mux21_comp_in_2(w_884), .mux21_comp_out(w_1125));
  mux21_comp #(.LEN(32))
    mux21_comp_1126 (.mux21_comp_sel(w_1120), .mux21_comp_in_1(w_1121), .mux21_comp_in_2(w_1125), .mux21_comp_out(w_1126));
  mux21_comp #(.LEN(32))
    mux21_comp_1127 (.mux21_comp_sel(w_1117), .mux21_comp_in_1(w_1118), .mux21_comp_in_2(w_1126), .mux21_comp_out(w_1127));
  mux21_comp #(.LEN(32))
    mux21_comp_1128 (.mux21_comp_sel(w_1114), .mux21_comp_in_1(w_1115), .mux21_comp_in_2(w_1127), .mux21_comp_out(w_1128));
  mux21_comp #(.LEN(32))
    mux21_comp_1129 (.mux21_comp_sel(w_1111), .mux21_comp_in_1(w_1112), .mux21_comp_in_2(w_1128), .mux21_comp_out(w_1129));
  mux21_comp #(.LEN(32))
    mux21_comp_1130 (.mux21_comp_sel(w_1108), .mux21_comp_in_1(w_1109), .mux21_comp_in_2(w_1129), .mux21_comp_out(w_1130));
  mux21_comp #(.LEN(32))
    mux21_comp_1131 (.mux21_comp_sel(w_1105), .mux21_comp_in_1(w_1106), .mux21_comp_in_2(w_1130), .mux21_comp_out(w_1131));
  mux21_comp #(.LEN(32))
    mux21_comp_1132 (.mux21_comp_sel(w_1102), .mux21_comp_in_1(w_1103), .mux21_comp_in_2(w_1131), .mux21_comp_out(w_1132));
  mux21_comp #(.LEN(32))
    mux21_comp_1133 (.mux21_comp_sel(w_1099), .mux21_comp_in_1(w_1100), .mux21_comp_in_2(w_1132), .mux21_comp_out(w_1133));
  mux21_comp #(.LEN(32))
    mux21_comp_1134 (.mux21_comp_sel(w_1096), .mux21_comp_in_1(w_1097), .mux21_comp_in_2(w_1133), .mux21_comp_out(w_1134));
  mux21_comp #(.LEN(32))
    mux21_comp_1135 (.mux21_comp_sel(w_1093), .mux21_comp_in_1(w_1094), .mux21_comp_in_2(w_1134), .mux21_comp_out(w_1135));
  mux21_comp #(.LEN(32))
    mux21_comp_1136 (.mux21_comp_sel(w_1090), .mux21_comp_in_1(w_1091), .mux21_comp_in_2(w_1135), .mux21_comp_out(w_1136));
  mux21_comp #(.LEN(32))
    mux21_comp_1137 (.mux21_comp_sel(w_1087), .mux21_comp_in_1(w_1088), .mux21_comp_in_2(w_1136), .mux21_comp_out(w_1137));
  mux21_comp #(.LEN(32))
    mux21_comp_1138 (.mux21_comp_sel(w_1084), .mux21_comp_in_1(w_1085), .mux21_comp_in_2(w_1137), .mux21_comp_out(w_1138));
  mux21_comp #(.LEN(32))
    mux21_comp_1139 (.mux21_comp_sel(w_1081), .mux21_comp_in_1(w_1082), .mux21_comp_in_2(w_1138), .mux21_comp_out(w_1139));
  mux21_comp #(.LEN(32))
    mux21_comp_1140 (.mux21_comp_sel(w_1078), .mux21_comp_in_1(w_1079), .mux21_comp_in_2(w_1139), .mux21_comp_out(w_1140));
  mux21_comp #(.LEN(32))
    mux21_comp_1141 (.mux21_comp_sel(w_1075), .mux21_comp_in_1(w_1076), .mux21_comp_in_2(w_1140), .mux21_comp_out(w_1141));
  mux21_comp #(.LEN(32))
    mux21_comp_1142 (.mux21_comp_sel(w_1072), .mux21_comp_in_1(w_1073), .mux21_comp_in_2(w_1141), .mux21_comp_out(w_1142));
  mux21_comp #(.LEN(32))
    mux21_comp_1143 (.mux21_comp_sel(w_1069), .mux21_comp_in_1(w_1070), .mux21_comp_in_2(w_1142), .mux21_comp_out(w_1143));
  mux21_comp #(.LEN(32))
    mux21_comp_1144 (.mux21_comp_sel(w_1066), .mux21_comp_in_1(w_1067), .mux21_comp_in_2(w_1143), .mux21_comp_out(w_1144));
  mux21_comp #(.LEN(32))
    mux21_comp_1145 (.mux21_comp_sel(w_1063), .mux21_comp_in_1(w_1064), .mux21_comp_in_2(w_1144), .mux21_comp_out(w_1145));
  mux21_comp #(.LEN(32))
    mux21_comp_1146 (.mux21_comp_sel(w_1060), .mux21_comp_in_1(w_1061), .mux21_comp_in_2(w_1145), .mux21_comp_out(w_1146));
  mux21_comp #(.LEN(32))
    mux21_comp_1147 (.mux21_comp_sel(w_1057), .mux21_comp_in_1(w_1058), .mux21_comp_in_2(w_1146), .mux21_comp_out(w_1147));
  mux21_comp #(.LEN(32))
    mux21_comp_1148 (.mux21_comp_sel(w_1054), .mux21_comp_in_1(w_1055), .mux21_comp_in_2(w_1147), .mux21_comp_out(w_1148));
  mux21_comp #(.LEN(32))
    mux21_comp_1149 (.mux21_comp_sel(w_1051), .mux21_comp_in_1(w_1052), .mux21_comp_in_2(w_1148), .mux21_comp_out(w_1149));
  mux21_comp #(.LEN(32))
    mux21_comp_1150 (.mux21_comp_sel(w_1048), .mux21_comp_in_1(w_1049), .mux21_comp_in_2(w_1149), .mux21_comp_out(w_1150));
  mux21_comp #(.LEN(32))
    mux21_comp_1151 (.mux21_comp_sel(w_1045), .mux21_comp_in_1(w_1046), .mux21_comp_in_2(w_1150), .mux21_comp_out(w_1151));
  mux21_comp #(.LEN(32))
    mux21_comp_1152 (.mux21_comp_sel(w_1042), .mux21_comp_in_1(w_1043), .mux21_comp_in_2(w_1151), .mux21_comp_out(w_1152));
  mux21_comp #(.LEN(32))
    mux21_comp_1153 (.mux21_comp_sel(w_1039), .mux21_comp_in_1(w_1040), .mux21_comp_in_2(w_1152), .mux21_comp_out(w_1153));
  mux21_comp #(.LEN(32))
    mux21_comp_1154 (.mux21_comp_sel(w_1036), .mux21_comp_in_1(w_1037), .mux21_comp_in_2(w_1153), .mux21_comp_out(w_1154));
  mux21_comp #(.LEN(32))
    mux21_comp_1155 (.mux21_comp_sel(w_1033), .mux21_comp_in_1(w_1034), .mux21_comp_in_2(w_1154), .mux21_comp_out(w_1155));
  slice #(.LEN(10), .LOWER(7), .UPPER(8))
    slice_1156 (.slice_in_1(w_883), .slice_out(w_1156));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1157 (.slice_in_1(w_885), .slice_out(w_1157));
  eq #(.LEN(5))
    eq_1158 (.eq_in_1(w_1157), .eq_in_2(5'd31), .eq_out(w_1158));
  sra #(.LEN(32), .SHAMT(31))
    sra_1159 (.sra_in_1(w_884), .sra_out(w_1159));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1160 (.slice_in_1(w_885), .slice_out(w_1160));
  eq #(.LEN(5))
    eq_1161 (.eq_in_1(w_1160), .eq_in_2(5'd30), .eq_out(w_1161));
  sra #(.LEN(32), .SHAMT(30))
    sra_1162 (.sra_in_1(w_884), .sra_out(w_1162));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1163 (.slice_in_1(w_885), .slice_out(w_1163));
  eq #(.LEN(5))
    eq_1164 (.eq_in_1(w_1163), .eq_in_2(5'd29), .eq_out(w_1164));
  sra #(.LEN(32), .SHAMT(29))
    sra_1165 (.sra_in_1(w_884), .sra_out(w_1165));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1166 (.slice_in_1(w_885), .slice_out(w_1166));
  eq #(.LEN(5))
    eq_1167 (.eq_in_1(w_1166), .eq_in_2(5'd28), .eq_out(w_1167));
  sra #(.LEN(32), .SHAMT(28))
    sra_1168 (.sra_in_1(w_884), .sra_out(w_1168));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1169 (.slice_in_1(w_885), .slice_out(w_1169));
  eq #(.LEN(5))
    eq_1170 (.eq_in_1(w_1169), .eq_in_2(5'd27), .eq_out(w_1170));
  sra #(.LEN(32), .SHAMT(27))
    sra_1171 (.sra_in_1(w_884), .sra_out(w_1171));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1172 (.slice_in_1(w_885), .slice_out(w_1172));
  eq #(.LEN(5))
    eq_1173 (.eq_in_1(w_1172), .eq_in_2(5'd26), .eq_out(w_1173));
  sra #(.LEN(32), .SHAMT(26))
    sra_1174 (.sra_in_1(w_884), .sra_out(w_1174));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1175 (.slice_in_1(w_885), .slice_out(w_1175));
  eq #(.LEN(5))
    eq_1176 (.eq_in_1(w_1175), .eq_in_2(5'd25), .eq_out(w_1176));
  sra #(.LEN(32), .SHAMT(25))
    sra_1177 (.sra_in_1(w_884), .sra_out(w_1177));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1178 (.slice_in_1(w_885), .slice_out(w_1178));
  eq #(.LEN(5))
    eq_1179 (.eq_in_1(w_1178), .eq_in_2(5'd24), .eq_out(w_1179));
  sra #(.LEN(32), .SHAMT(24))
    sra_1180 (.sra_in_1(w_884), .sra_out(w_1180));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1181 (.slice_in_1(w_885), .slice_out(w_1181));
  eq #(.LEN(5))
    eq_1182 (.eq_in_1(w_1181), .eq_in_2(5'd23), .eq_out(w_1182));
  sra #(.LEN(32), .SHAMT(23))
    sra_1183 (.sra_in_1(w_884), .sra_out(w_1183));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1184 (.slice_in_1(w_885), .slice_out(w_1184));
  eq #(.LEN(5))
    eq_1185 (.eq_in_1(w_1184), .eq_in_2(5'd22), .eq_out(w_1185));
  sra #(.LEN(32), .SHAMT(22))
    sra_1186 (.sra_in_1(w_884), .sra_out(w_1186));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1187 (.slice_in_1(w_885), .slice_out(w_1187));
  eq #(.LEN(5))
    eq_1188 (.eq_in_1(w_1187), .eq_in_2(5'd21), .eq_out(w_1188));
  sra #(.LEN(32), .SHAMT(21))
    sra_1189 (.sra_in_1(w_884), .sra_out(w_1189));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1190 (.slice_in_1(w_885), .slice_out(w_1190));
  eq #(.LEN(5))
    eq_1191 (.eq_in_1(w_1190), .eq_in_2(5'd20), .eq_out(w_1191));
  sra #(.LEN(32), .SHAMT(20))
    sra_1192 (.sra_in_1(w_884), .sra_out(w_1192));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1193 (.slice_in_1(w_885), .slice_out(w_1193));
  eq #(.LEN(5))
    eq_1194 (.eq_in_1(w_1193), .eq_in_2(5'd19), .eq_out(w_1194));
  sra #(.LEN(32), .SHAMT(19))
    sra_1195 (.sra_in_1(w_884), .sra_out(w_1195));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1196 (.slice_in_1(w_885), .slice_out(w_1196));
  eq #(.LEN(5))
    eq_1197 (.eq_in_1(w_1196), .eq_in_2(5'd18), .eq_out(w_1197));
  sra #(.LEN(32), .SHAMT(18))
    sra_1198 (.sra_in_1(w_884), .sra_out(w_1198));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1199 (.slice_in_1(w_885), .slice_out(w_1199));
  eq #(.LEN(5))
    eq_1200 (.eq_in_1(w_1199), .eq_in_2(5'd17), .eq_out(w_1200));
  sra #(.LEN(32), .SHAMT(17))
    sra_1201 (.sra_in_1(w_884), .sra_out(w_1201));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1202 (.slice_in_1(w_885), .slice_out(w_1202));
  eq #(.LEN(5))
    eq_1203 (.eq_in_1(w_1202), .eq_in_2(5'd16), .eq_out(w_1203));
  sra #(.LEN(32), .SHAMT(16))
    sra_1204 (.sra_in_1(w_884), .sra_out(w_1204));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1205 (.slice_in_1(w_885), .slice_out(w_1205));
  eq #(.LEN(5))
    eq_1206 (.eq_in_1(w_1205), .eq_in_2(5'd15), .eq_out(w_1206));
  sra #(.LEN(32), .SHAMT(15))
    sra_1207 (.sra_in_1(w_884), .sra_out(w_1207));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1208 (.slice_in_1(w_885), .slice_out(w_1208));
  eq #(.LEN(5))
    eq_1209 (.eq_in_1(w_1208), .eq_in_2(5'd14), .eq_out(w_1209));
  sra #(.LEN(32), .SHAMT(14))
    sra_1210 (.sra_in_1(w_884), .sra_out(w_1210));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1211 (.slice_in_1(w_885), .slice_out(w_1211));
  eq #(.LEN(5))
    eq_1212 (.eq_in_1(w_1211), .eq_in_2(5'd13), .eq_out(w_1212));
  sra #(.LEN(32), .SHAMT(13))
    sra_1213 (.sra_in_1(w_884), .sra_out(w_1213));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1214 (.slice_in_1(w_885), .slice_out(w_1214));
  eq #(.LEN(5))
    eq_1215 (.eq_in_1(w_1214), .eq_in_2(5'd12), .eq_out(w_1215));
  sra #(.LEN(32), .SHAMT(12))
    sra_1216 (.sra_in_1(w_884), .sra_out(w_1216));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1217 (.slice_in_1(w_885), .slice_out(w_1217));
  eq #(.LEN(5))
    eq_1218 (.eq_in_1(w_1217), .eq_in_2(5'd11), .eq_out(w_1218));
  sra #(.LEN(32), .SHAMT(11))
    sra_1219 (.sra_in_1(w_884), .sra_out(w_1219));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1220 (.slice_in_1(w_885), .slice_out(w_1220));
  eq #(.LEN(5))
    eq_1221 (.eq_in_1(w_1220), .eq_in_2(5'd10), .eq_out(w_1221));
  sra #(.LEN(32), .SHAMT(10))
    sra_1222 (.sra_in_1(w_884), .sra_out(w_1222));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1223 (.slice_in_1(w_885), .slice_out(w_1223));
  eq #(.LEN(5))
    eq_1224 (.eq_in_1(w_1223), .eq_in_2(5'd9), .eq_out(w_1224));
  sra #(.LEN(32), .SHAMT(9))
    sra_1225 (.sra_in_1(w_884), .sra_out(w_1225));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1226 (.slice_in_1(w_885), .slice_out(w_1226));
  eq #(.LEN(5))
    eq_1227 (.eq_in_1(w_1226), .eq_in_2(5'd8), .eq_out(w_1227));
  sra #(.LEN(32), .SHAMT(8))
    sra_1228 (.sra_in_1(w_884), .sra_out(w_1228));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1229 (.slice_in_1(w_885), .slice_out(w_1229));
  eq #(.LEN(5))
    eq_1230 (.eq_in_1(w_1229), .eq_in_2(5'd7), .eq_out(w_1230));
  sra #(.LEN(32), .SHAMT(7))
    sra_1231 (.sra_in_1(w_884), .sra_out(w_1231));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1232 (.slice_in_1(w_885), .slice_out(w_1232));
  eq #(.LEN(5))
    eq_1233 (.eq_in_1(w_1232), .eq_in_2(5'd6), .eq_out(w_1233));
  sra #(.LEN(32), .SHAMT(6))
    sra_1234 (.sra_in_1(w_884), .sra_out(w_1234));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1235 (.slice_in_1(w_885), .slice_out(w_1235));
  eq #(.LEN(5))
    eq_1236 (.eq_in_1(w_1235), .eq_in_2(5'd5), .eq_out(w_1236));
  sra #(.LEN(32), .SHAMT(5))
    sra_1237 (.sra_in_1(w_884), .sra_out(w_1237));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1238 (.slice_in_1(w_885), .slice_out(w_1238));
  eq #(.LEN(5))
    eq_1239 (.eq_in_1(w_1238), .eq_in_2(5'd4), .eq_out(w_1239));
  sra #(.LEN(32), .SHAMT(4))
    sra_1240 (.sra_in_1(w_884), .sra_out(w_1240));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1241 (.slice_in_1(w_885), .slice_out(w_1241));
  eq #(.LEN(5))
    eq_1242 (.eq_in_1(w_1241), .eq_in_2(5'd3), .eq_out(w_1242));
  sra #(.LEN(32), .SHAMT(3))
    sra_1243 (.sra_in_1(w_884), .sra_out(w_1243));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1244 (.slice_in_1(w_885), .slice_out(w_1244));
  eq #(.LEN(5))
    eq_1245 (.eq_in_1(w_1244), .eq_in_2(5'd2), .eq_out(w_1245));
  sra #(.LEN(32), .SHAMT(2))
    sra_1246 (.sra_in_1(w_884), .sra_out(w_1246));
  slice #(.LEN(32), .LOWER(0), .UPPER(5))
    slice_1247 (.slice_in_1(w_885), .slice_out(w_1247));
  eq #(.LEN(5))
    eq_1248 (.eq_in_1(w_1247), .eq_in_2(5'd1), .eq_out(w_1248));
  sra #(.LEN(32), .SHAMT(1))
    sra_1249 (.sra_in_1(w_884), .sra_out(w_1249));
  mux21_comp #(.LEN(32))
    mux21_comp_1250 (.mux21_comp_sel(w_1248), .mux21_comp_in_1(w_1249), .mux21_comp_in_2(w_884), .mux21_comp_out(w_1250));
  mux21_comp #(.LEN(32))
    mux21_comp_1251 (.mux21_comp_sel(w_1245), .mux21_comp_in_1(w_1246), .mux21_comp_in_2(w_1250), .mux21_comp_out(w_1251));
  mux21_comp #(.LEN(32))
    mux21_comp_1252 (.mux21_comp_sel(w_1242), .mux21_comp_in_1(w_1243), .mux21_comp_in_2(w_1251), .mux21_comp_out(w_1252));
  mux21_comp #(.LEN(32))
    mux21_comp_1253 (.mux21_comp_sel(w_1239), .mux21_comp_in_1(w_1240), .mux21_comp_in_2(w_1252), .mux21_comp_out(w_1253));
  mux21_comp #(.LEN(32))
    mux21_comp_1254 (.mux21_comp_sel(w_1236), .mux21_comp_in_1(w_1237), .mux21_comp_in_2(w_1253), .mux21_comp_out(w_1254));
  mux21_comp #(.LEN(32))
    mux21_comp_1255 (.mux21_comp_sel(w_1233), .mux21_comp_in_1(w_1234), .mux21_comp_in_2(w_1254), .mux21_comp_out(w_1255));
  mux21_comp #(.LEN(32))
    mux21_comp_1256 (.mux21_comp_sel(w_1230), .mux21_comp_in_1(w_1231), .mux21_comp_in_2(w_1255), .mux21_comp_out(w_1256));
  mux21_comp #(.LEN(32))
    mux21_comp_1257 (.mux21_comp_sel(w_1227), .mux21_comp_in_1(w_1228), .mux21_comp_in_2(w_1256), .mux21_comp_out(w_1257));
  mux21_comp #(.LEN(32))
    mux21_comp_1258 (.mux21_comp_sel(w_1224), .mux21_comp_in_1(w_1225), .mux21_comp_in_2(w_1257), .mux21_comp_out(w_1258));
  mux21_comp #(.LEN(32))
    mux21_comp_1259 (.mux21_comp_sel(w_1221), .mux21_comp_in_1(w_1222), .mux21_comp_in_2(w_1258), .mux21_comp_out(w_1259));
  mux21_comp #(.LEN(32))
    mux21_comp_1260 (.mux21_comp_sel(w_1218), .mux21_comp_in_1(w_1219), .mux21_comp_in_2(w_1259), .mux21_comp_out(w_1260));
  mux21_comp #(.LEN(32))
    mux21_comp_1261 (.mux21_comp_sel(w_1215), .mux21_comp_in_1(w_1216), .mux21_comp_in_2(w_1260), .mux21_comp_out(w_1261));
  mux21_comp #(.LEN(32))
    mux21_comp_1262 (.mux21_comp_sel(w_1212), .mux21_comp_in_1(w_1213), .mux21_comp_in_2(w_1261), .mux21_comp_out(w_1262));
  mux21_comp #(.LEN(32))
    mux21_comp_1263 (.mux21_comp_sel(w_1209), .mux21_comp_in_1(w_1210), .mux21_comp_in_2(w_1262), .mux21_comp_out(w_1263));
  mux21_comp #(.LEN(32))
    mux21_comp_1264 (.mux21_comp_sel(w_1206), .mux21_comp_in_1(w_1207), .mux21_comp_in_2(w_1263), .mux21_comp_out(w_1264));
  mux21_comp #(.LEN(32))
    mux21_comp_1265 (.mux21_comp_sel(w_1203), .mux21_comp_in_1(w_1204), .mux21_comp_in_2(w_1264), .mux21_comp_out(w_1265));
  mux21_comp #(.LEN(32))
    mux21_comp_1266 (.mux21_comp_sel(w_1200), .mux21_comp_in_1(w_1201), .mux21_comp_in_2(w_1265), .mux21_comp_out(w_1266));
  mux21_comp #(.LEN(32))
    mux21_comp_1267 (.mux21_comp_sel(w_1197), .mux21_comp_in_1(w_1198), .mux21_comp_in_2(w_1266), .mux21_comp_out(w_1267));
  mux21_comp #(.LEN(32))
    mux21_comp_1268 (.mux21_comp_sel(w_1194), .mux21_comp_in_1(w_1195), .mux21_comp_in_2(w_1267), .mux21_comp_out(w_1268));
  mux21_comp #(.LEN(32))
    mux21_comp_1269 (.mux21_comp_sel(w_1191), .mux21_comp_in_1(w_1192), .mux21_comp_in_2(w_1268), .mux21_comp_out(w_1269));
  mux21_comp #(.LEN(32))
    mux21_comp_1270 (.mux21_comp_sel(w_1188), .mux21_comp_in_1(w_1189), .mux21_comp_in_2(w_1269), .mux21_comp_out(w_1270));
  mux21_comp #(.LEN(32))
    mux21_comp_1271 (.mux21_comp_sel(w_1185), .mux21_comp_in_1(w_1186), .mux21_comp_in_2(w_1270), .mux21_comp_out(w_1271));
  mux21_comp #(.LEN(32))
    mux21_comp_1272 (.mux21_comp_sel(w_1182), .mux21_comp_in_1(w_1183), .mux21_comp_in_2(w_1271), .mux21_comp_out(w_1272));
  mux21_comp #(.LEN(32))
    mux21_comp_1273 (.mux21_comp_sel(w_1179), .mux21_comp_in_1(w_1180), .mux21_comp_in_2(w_1272), .mux21_comp_out(w_1273));
  mux21_comp #(.LEN(32))
    mux21_comp_1274 (.mux21_comp_sel(w_1176), .mux21_comp_in_1(w_1177), .mux21_comp_in_2(w_1273), .mux21_comp_out(w_1274));
  mux21_comp #(.LEN(32))
    mux21_comp_1275 (.mux21_comp_sel(w_1173), .mux21_comp_in_1(w_1174), .mux21_comp_in_2(w_1274), .mux21_comp_out(w_1275));
  mux21_comp #(.LEN(32))
    mux21_comp_1276 (.mux21_comp_sel(w_1170), .mux21_comp_in_1(w_1171), .mux21_comp_in_2(w_1275), .mux21_comp_out(w_1276));
  mux21_comp #(.LEN(32))
    mux21_comp_1277 (.mux21_comp_sel(w_1167), .mux21_comp_in_1(w_1168), .mux21_comp_in_2(w_1276), .mux21_comp_out(w_1277));
  mux21_comp #(.LEN(32))
    mux21_comp_1278 (.mux21_comp_sel(w_1164), .mux21_comp_in_1(w_1165), .mux21_comp_in_2(w_1277), .mux21_comp_out(w_1278));
  mux21_comp #(.LEN(32))
    mux21_comp_1279 (.mux21_comp_sel(w_1161), .mux21_comp_in_1(w_1162), .mux21_comp_in_2(w_1278), .mux21_comp_out(w_1279));
  mux21_comp #(.LEN(32))
    mux21_comp_1280 (.mux21_comp_sel(w_1158), .mux21_comp_in_1(w_1159), .mux21_comp_in_2(w_1279), .mux21_comp_out(w_1280));
  slice #(.LEN(10), .LOWER(8), .UPPER(9))
    slice_1281 (.slice_in_1(w_883), .slice_out(w_1281));
  or_comp #(.LEN(32))
    or_comp_1282 (.or_comp_in_1(w_884), .or_comp_in_2(w_885), .or_comp_out(w_1282));
  and_comp #(.LEN(32))
    and_comp_1283 (.and_comp_in_1(w_884), .and_comp_in_2(w_885), .and_comp_out(w_1283));
  mux21_comp #(.LEN(32))
    mux21_comp_1284 (.mux21_comp_sel(w_1281), .mux21_comp_in_1(w_1282), .mux21_comp_in_2(w_1283), .mux21_comp_out(w_1284));
  mux21_comp #(.LEN(32))
    mux21_comp_1285 (.mux21_comp_sel(w_1156), .mux21_comp_in_1(w_1280), .mux21_comp_in_2(w_1284), .mux21_comp_out(w_1285));
  mux21_comp #(.LEN(32))
    mux21_comp_1286 (.mux21_comp_sel(w_1031), .mux21_comp_in_1(w_1155), .mux21_comp_in_2(w_1285), .mux21_comp_out(w_1286));
  mux21_comp #(.LEN(32))
    mux21_comp_1287 (.mux21_comp_sel(w_906), .mux21_comp_in_1(w_1030), .mux21_comp_in_2(w_1286), .mux21_comp_out(w_1287));
  mux21_comp #(.LEN(32))
    mux21_comp_1288 (.mux21_comp_sel(w_904), .mux21_comp_in_1(w_905), .mux21_comp_in_2(w_1287), .mux21_comp_out(w_1288));
  mux21_comp #(.LEN(32))
    mux21_comp_1289 (.mux21_comp_sel(w_901), .mux21_comp_in_1(w_903), .mux21_comp_in_2(w_1288), .mux21_comp_out(w_1289));
  mux21_comp #(.LEN(32))
    mux21_comp_1290 (.mux21_comp_sel(w_898), .mux21_comp_in_1(w_900), .mux21_comp_in_2(w_1289), .mux21_comp_out(w_1290));
  mux21_comp #(.LEN(32))
    mux21_comp_1291 (.mux21_comp_sel(w_890), .mux21_comp_in_1(w_897), .mux21_comp_in_2(w_1290), .mux21_comp_out(w_1291));
  mux21_comp #(.LEN(32))
    mux21_comp_1292 (.mux21_comp_sel(w_886), .mux21_comp_in_1(w_889), .mux21_comp_in_2(w_1291), .mux21_comp_out(w_1292));
  mux21_comp #(.LEN(32))
    mux21_comp_1293 (.mux21_comp_sel(w_849), .mux21_comp_in_1(w_1292), .mux21_comp_in_2(32'd0), .mux21_comp_out(w_1293));
  mux21_comp #(.LEN(32))
    mux21_comp_1294 (.mux21_comp_sel(w_841), .mux21_comp_in_1(w_844), .mux21_comp_in_2(w_1293), .mux21_comp_out(w_1294));
  mux21_comp #(.LEN(32))
    mux21_comp_1295 (.mux21_comp_sel(w_833), .mux21_comp_in_1(w_836), .mux21_comp_in_2(w_1294), .mux21_comp_out(w_1295));
  mux21_comp #(.LEN(32))
    mux21_comp_1296 (.mux21_comp_sel(w_831), .mux21_comp_in_1(w_595), .mux21_comp_in_2(w_1295), .mux21_comp_out(w_1296));
  mux21_comp #(.LEN(32))
    mux21_comp_1297 (.mux21_comp_sel(w_473), .mux21_comp_in_1(w_829), .mux21_comp_in_2(w_1296), .mux21_comp_out(w_1297));
  not_comp #(.LEN(1))
    not_comp_1298 (.not_comp_in_1(w_0), .not_comp_out(w_1298));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_1299 (.slice_in_1(w_1), .slice_out(w_1299));
  eq #(.LEN(7))
    eq_1300 (.eq_in_1(w_1299), .eq_in_2(7'd35), .eq_out(w_1300));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_1301 (.slice_in_1(w_1), .slice_out(w_1301));
  eq #(.LEN(7))
    eq_1302 (.eq_in_1(w_1301), .eq_in_2(7'd3), .eq_out(w_1302));
  or_comp #(.LEN(1))
    or_comp_1303 (.or_comp_in_1(w_1300), .or_comp_in_2(w_1302), .or_comp_out(w_1303));
  mux21_comp #(.LEN(1))
    mux21_comp_1304 (.mux21_comp_sel(w_1303), .mux21_comp_in_1(1'd1), .mux21_comp_in_2(1'd0), .mux21_comp_out(w_1304));
  mux21_comp #(.LEN(1))
    mux21_comp_1305 (.mux21_comp_sel(w_473), .mux21_comp_in_1(1'd0), .mux21_comp_in_2(w_1304), .mux21_comp_out(w_1305));
  mux21_comp #(.LEN(1))
    mux21_comp_1306 (.mux21_comp_sel(w_1298), .mux21_comp_in_1(1'd0), .mux21_comp_in_2(w_1305), .mux21_comp_out(w_1306));
  not_comp #(.LEN(1))
    not_comp_1307 (.not_comp_in_1(w_0), .not_comp_out(w_1307));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_1308 (.slice_in_1(w_1), .slice_out(w_1308));
  eq #(.LEN(7))
    eq_1309 (.eq_in_1(w_1308), .eq_in_2(7'd35), .eq_out(w_1309));
  mux21_comp #(.LEN(1))
    mux21_comp_1310 (.mux21_comp_sel(w_1309), .mux21_comp_in_1(1'd1), .mux21_comp_in_2(1'd0), .mux21_comp_out(w_1310));
  mux21_comp #(.LEN(1))
    mux21_comp_1311 (.mux21_comp_sel(w_473), .mux21_comp_in_1(1'd0), .mux21_comp_in_2(w_1310), .mux21_comp_out(w_1311));
  mux21_comp #(.LEN(1))
    mux21_comp_1312 (.mux21_comp_sel(w_1307), .mux21_comp_in_1(1'd0), .mux21_comp_in_2(w_1311), .mux21_comp_out(w_1312));
  not_comp #(.LEN(1))
    not_comp_1313 (.not_comp_in_1(w_0), .not_comp_out(w_1313));
  slice #(.LEN(32), .LOWER(0), .UPPER(7))
    slice_1314 (.slice_in_1(w_1), .slice_out(w_1314));
  eq #(.LEN(7))
    eq_1315 (.eq_in_1(w_1314), .eq_in_2(7'd35), .eq_out(w_1315));
  slice #(.LEN(32), .LOWER(20), .UPPER(25))
    slice_1316 (.slice_in_1(w_1), .slice_out(w_1316));
  slice #(.LEN(32), .LOWER(7), .UPPER(12))
    slice_1317 (.slice_in_1(w_1), .slice_out(w_1317));
  mux21_comp #(.LEN(5))
    mux21_comp_1318 (.mux21_comp_sel(w_1315), .mux21_comp_in_1(w_1316), .mux21_comp_in_2(w_1317), .mux21_comp_out(w_1318));
  mux21_comp #(.LEN(5))
    mux21_comp_1319 (.mux21_comp_sel(w_1313), .mux21_comp_in_1(5'd0), .mux21_comp_in_2(w_1318), .mux21_comp_out(w_1319));
  not_comp #(.LEN(1))
    not_comp_1320 (.not_comp_in_1(w_0), .not_comp_out(w_1320));
  mux21_comp #(.LEN(32))
    mux21_comp_1321 (.mux21_comp_sel(w_1320), .mux21_comp_in_1(32'd0), .mux21_comp_in_2(w_472), .mux21_comp_out(w_1321));
  not_comp #(.LEN(1))
    not_comp_1322 (.not_comp_in_1(w_0), .not_comp_out(w_1322));
  add #(.LEN(32))
    add_1323 (.add_in_1(w_2), .add_in_2(32'd4), .add_out(w_1323));
  slice #(.LEN(33), .LOWER(0), .UPPER(32))
    slice_1325 (.slice_in_1(w_1324), .slice_out(w_1325));
  mux21_comp #(.LEN(32))
    mux21_comp_1326 (.mux21_comp_sel(w_1322), .mux21_comp_in_1(32'd0), .mux21_comp_in_2(w_1325), .mux21_comp_out(w_1326));
  not_comp #(.LEN(1))
    not_comp_1327 (.not_comp_in_1(w_0), .not_comp_out(w_1327));
  slice #(.LEN(32), .LOWER(12), .UPPER(15))
    slice_1328 (.slice_in_1(w_1), .slice_out(w_1328));
  mux21_comp #(.LEN(3))
    mux21_comp_1329 (.mux21_comp_sel(w_1327), .mux21_comp_in_1(3'd0), .mux21_comp_in_2(w_1328), .mux21_comp_out(w_1329));
  eq #(.LEN(5))
    eq_1452 (.eq_in_1(w_1386), .eq_in_2(5'd31), .eq_out(w_1452));
  mux21_comp #(.LEN(32))
    mux21_comp_1453 (.mux21_comp_sel(w_1452), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1420), .mux21_comp_out(w_1453));
  eq #(.LEN(5))
    eq_1454 (.eq_in_1(w_1386), .eq_in_2(5'd30), .eq_out(w_1454));
  mux21_comp #(.LEN(32))
    mux21_comp_1455 (.mux21_comp_sel(w_1454), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1421), .mux21_comp_out(w_1455));
  eq #(.LEN(5))
    eq_1456 (.eq_in_1(w_1386), .eq_in_2(5'd29), .eq_out(w_1456));
  mux21_comp #(.LEN(32))
    mux21_comp_1457 (.mux21_comp_sel(w_1456), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1422), .mux21_comp_out(w_1457));
  eq #(.LEN(5))
    eq_1458 (.eq_in_1(w_1386), .eq_in_2(5'd28), .eq_out(w_1458));
  mux21_comp #(.LEN(32))
    mux21_comp_1459 (.mux21_comp_sel(w_1458), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1423), .mux21_comp_out(w_1459));
  eq #(.LEN(5))
    eq_1460 (.eq_in_1(w_1386), .eq_in_2(5'd27), .eq_out(w_1460));
  mux21_comp #(.LEN(32))
    mux21_comp_1461 (.mux21_comp_sel(w_1460), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1424), .mux21_comp_out(w_1461));
  eq #(.LEN(5))
    eq_1462 (.eq_in_1(w_1386), .eq_in_2(5'd26), .eq_out(w_1462));
  mux21_comp #(.LEN(32))
    mux21_comp_1463 (.mux21_comp_sel(w_1462), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1425), .mux21_comp_out(w_1463));
  eq #(.LEN(5))
    eq_1464 (.eq_in_1(w_1386), .eq_in_2(5'd25), .eq_out(w_1464));
  mux21_comp #(.LEN(32))
    mux21_comp_1465 (.mux21_comp_sel(w_1464), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1426), .mux21_comp_out(w_1465));
  eq #(.LEN(5))
    eq_1466 (.eq_in_1(w_1386), .eq_in_2(5'd24), .eq_out(w_1466));
  mux21_comp #(.LEN(32))
    mux21_comp_1467 (.mux21_comp_sel(w_1466), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1427), .mux21_comp_out(w_1467));
  eq #(.LEN(5))
    eq_1468 (.eq_in_1(w_1386), .eq_in_2(5'd23), .eq_out(w_1468));
  mux21_comp #(.LEN(32))
    mux21_comp_1469 (.mux21_comp_sel(w_1468), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1428), .mux21_comp_out(w_1469));
  eq #(.LEN(5))
    eq_1470 (.eq_in_1(w_1386), .eq_in_2(5'd22), .eq_out(w_1470));
  mux21_comp #(.LEN(32))
    mux21_comp_1471 (.mux21_comp_sel(w_1470), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1429), .mux21_comp_out(w_1471));
  eq #(.LEN(5))
    eq_1472 (.eq_in_1(w_1386), .eq_in_2(5'd21), .eq_out(w_1472));
  mux21_comp #(.LEN(32))
    mux21_comp_1473 (.mux21_comp_sel(w_1472), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1430), .mux21_comp_out(w_1473));
  eq #(.LEN(5))
    eq_1474 (.eq_in_1(w_1386), .eq_in_2(5'd20), .eq_out(w_1474));
  mux21_comp #(.LEN(32))
    mux21_comp_1475 (.mux21_comp_sel(w_1474), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1431), .mux21_comp_out(w_1475));
  eq #(.LEN(5))
    eq_1476 (.eq_in_1(w_1386), .eq_in_2(5'd19), .eq_out(w_1476));
  mux21_comp #(.LEN(32))
    mux21_comp_1477 (.mux21_comp_sel(w_1476), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1432), .mux21_comp_out(w_1477));
  eq #(.LEN(5))
    eq_1478 (.eq_in_1(w_1386), .eq_in_2(5'd18), .eq_out(w_1478));
  mux21_comp #(.LEN(32))
    mux21_comp_1479 (.mux21_comp_sel(w_1478), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1433), .mux21_comp_out(w_1479));
  eq #(.LEN(5))
    eq_1480 (.eq_in_1(w_1386), .eq_in_2(5'd17), .eq_out(w_1480));
  mux21_comp #(.LEN(32))
    mux21_comp_1481 (.mux21_comp_sel(w_1480), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1434), .mux21_comp_out(w_1481));
  eq #(.LEN(5))
    eq_1482 (.eq_in_1(w_1386), .eq_in_2(5'd16), .eq_out(w_1482));
  mux21_comp #(.LEN(32))
    mux21_comp_1483 (.mux21_comp_sel(w_1482), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1435), .mux21_comp_out(w_1483));
  eq #(.LEN(5))
    eq_1484 (.eq_in_1(w_1386), .eq_in_2(5'd15), .eq_out(w_1484));
  mux21_comp #(.LEN(32))
    mux21_comp_1485 (.mux21_comp_sel(w_1484), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1436), .mux21_comp_out(w_1485));
  eq #(.LEN(5))
    eq_1486 (.eq_in_1(w_1386), .eq_in_2(5'd14), .eq_out(w_1486));
  mux21_comp #(.LEN(32))
    mux21_comp_1487 (.mux21_comp_sel(w_1486), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1437), .mux21_comp_out(w_1487));
  eq #(.LEN(5))
    eq_1488 (.eq_in_1(w_1386), .eq_in_2(5'd13), .eq_out(w_1488));
  mux21_comp #(.LEN(32))
    mux21_comp_1489 (.mux21_comp_sel(w_1488), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1438), .mux21_comp_out(w_1489));
  eq #(.LEN(5))
    eq_1490 (.eq_in_1(w_1386), .eq_in_2(5'd12), .eq_out(w_1490));
  mux21_comp #(.LEN(32))
    mux21_comp_1491 (.mux21_comp_sel(w_1490), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1439), .mux21_comp_out(w_1491));
  eq #(.LEN(5))
    eq_1492 (.eq_in_1(w_1386), .eq_in_2(5'd11), .eq_out(w_1492));
  mux21_comp #(.LEN(32))
    mux21_comp_1493 (.mux21_comp_sel(w_1492), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1440), .mux21_comp_out(w_1493));
  eq #(.LEN(5))
    eq_1494 (.eq_in_1(w_1386), .eq_in_2(5'd10), .eq_out(w_1494));
  mux21_comp #(.LEN(32))
    mux21_comp_1495 (.mux21_comp_sel(w_1494), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1441), .mux21_comp_out(w_1495));
  eq #(.LEN(5))
    eq_1496 (.eq_in_1(w_1386), .eq_in_2(5'd9), .eq_out(w_1496));
  mux21_comp #(.LEN(32))
    mux21_comp_1497 (.mux21_comp_sel(w_1496), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1442), .mux21_comp_out(w_1497));
  eq #(.LEN(5))
    eq_1498 (.eq_in_1(w_1386), .eq_in_2(5'd8), .eq_out(w_1498));
  mux21_comp #(.LEN(32))
    mux21_comp_1499 (.mux21_comp_sel(w_1498), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1443), .mux21_comp_out(w_1499));
  eq #(.LEN(5))
    eq_1500 (.eq_in_1(w_1386), .eq_in_2(5'd7), .eq_out(w_1500));
  mux21_comp #(.LEN(32))
    mux21_comp_1501 (.mux21_comp_sel(w_1500), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1444), .mux21_comp_out(w_1501));
  eq #(.LEN(5))
    eq_1502 (.eq_in_1(w_1386), .eq_in_2(5'd6), .eq_out(w_1502));
  mux21_comp #(.LEN(32))
    mux21_comp_1503 (.mux21_comp_sel(w_1502), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1445), .mux21_comp_out(w_1503));
  eq #(.LEN(5))
    eq_1504 (.eq_in_1(w_1386), .eq_in_2(5'd5), .eq_out(w_1504));
  mux21_comp #(.LEN(32))
    mux21_comp_1505 (.mux21_comp_sel(w_1504), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1446), .mux21_comp_out(w_1505));
  eq #(.LEN(5))
    eq_1506 (.eq_in_1(w_1386), .eq_in_2(5'd4), .eq_out(w_1506));
  mux21_comp #(.LEN(32))
    mux21_comp_1507 (.mux21_comp_sel(w_1506), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1447), .mux21_comp_out(w_1507));
  eq #(.LEN(5))
    eq_1508 (.eq_in_1(w_1386), .eq_in_2(5'd3), .eq_out(w_1508));
  mux21_comp #(.LEN(32))
    mux21_comp_1509 (.mux21_comp_sel(w_1508), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1448), .mux21_comp_out(w_1509));
  eq #(.LEN(5))
    eq_1510 (.eq_in_1(w_1386), .eq_in_2(5'd2), .eq_out(w_1510));
  mux21_comp #(.LEN(32))
    mux21_comp_1511 (.mux21_comp_sel(w_1510), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1449), .mux21_comp_out(w_1511));
  eq #(.LEN(5))
    eq_1512 (.eq_in_1(w_1386), .eq_in_2(5'd1), .eq_out(w_1512));
  mux21_comp #(.LEN(32))
    mux21_comp_1513 (.mux21_comp_sel(w_1512), .mux21_comp_in_1(w_1387), .mux21_comp_in_2(w_1450), .mux21_comp_out(w_1513));

  always @ (posedge clk) begin
    r_3 <= w_1579;
    r_4 <= w_1580;
    r_5 <= w_1581;
    r_6 <= w_1582;
    r_7 <= w_1583;
    r_8 <= w_1584;
    r_9 <= w_1585;
    r_10 <= w_1586;
    r_11 <= w_1587;
    r_12 <= w_1588;
    r_13 <= w_1589;
    r_14 <= w_1590;
    r_15 <= w_1591;
    r_16 <= w_1592;
    r_17 <= w_1593;
    r_18 <= w_1594;
    r_19 <= w_1595;
    r_20 <= w_1596;
    r_21 <= w_1597;
    r_22 <= w_1598;
    r_23 <= w_1599;
    r_24 <= w_1600;
    r_25 <= w_1601;
    r_26 <= w_1602;
    r_27 <= w_1603;
    r_28 <= w_1604;
    r_29 <= w_1605;
    r_30 <= w_1606;
    r_31 <= w_1607;
    r_32 <= w_1608;
    r_33 <= w_1609;
    r_34 <= w_1610;
    r_459 <= w_1620;
    r_460 <= w_1621;
    r_461 <= w_1622;
    r_462 <= w_1623;
    r_463 <= w_1624;
    r_464 <= w_1625;
end

endmodule
